	// verilator_coverage annotation
	module ALU( // @[:@3.2]
%000002	  input  [5:0]  io_opcode, // @[:@6.4]
%000060	  input  [63:0] io_in1, // @[:@6.4]
%000060	  input  [63:0] io_in2, // @[:@6.4]
%000062	  output [63:0] io_out, // @[:@6.4]
%000003	  output        io_zero // @[:@6.4]
	);
	  wire  _T_15; // @[ALUop.scala 20:29:@8.4]
	  wire [63:0] _T_16; // @[ALU.scala 19:54:@9.4]
	  wire [64:0] _T_18; // @[ALU.scala 19:62:@10.4]
	  wire [63:0] _T_19; // @[ALU.scala 19:62:@11.4]
	  wire [63:0] _T_20; // @[ALU.scala 19:35:@12.4]
%000062	  wire [64:0] add_result; // @[ALU.scala 19:29:@13.4]
%000060	  wire [63:0] xor_result; // @[ALU.scala 20:29:@14.4]
%000060	  wire [63:0] or_result; // @[ALU.scala 21:29:@15.4]
%000060	  wire [63:0] and_result; // @[ALU.scala 22:29:@16.4]
	  wire  _T_21; // @[ALU.scala 24:41:@17.4]
%000001	  wire  sltu_result; // @[ALU.scala 24:30:@18.4]
	  wire  _T_22; // @[ALU.scala 25:40:@19.4]
%000001	  wire  slt_result; // @[ALU.scala 25:51:@20.4]
%000006	  wire [4:0] shamt; // @[ALU.scala 28:23:@21.4]
	  wire [94:0] _GEN_0; // @[ALU.scala 29:30:@22.4]
	  wire [94:0] _T_23; // @[ALU.scala 29:30:@22.4]
%000060	  wire [63:0] sll_result; // @[ALU.scala 29:39:@23.4]
	  wire [63:0] _T_24; // @[ALU.scala 30:36:@24.4]
	  wire [63:0] _T_25; // @[ALU.scala 30:39:@25.4]
%000008	  wire [63:0] sra_result; // @[ALU.scala 30:55:@26.4]
%000008	  wire [63:0] srl_result; // @[ALU.scala 31:29:@27.4]
	  wire [63:0] _T_26; // @[ALU.scala 33:33:@28.4]
	  wire  _T_28; // @[ALU.scala 34:20:@29.4]
	  wire [63:0] _T_30; // @[Cat.scala 30:58:@30.4]
	  wire  _T_32; // @[ALU.scala 35:20:@31.4]
	  wire [63:0] _T_34; // @[Cat.scala 30:58:@32.4]
	  wire  _T_36; // @[ALU.scala 36:20:@33.4]
	  wire  _T_38; // @[ALU.scala 37:20:@34.4]
	  wire  _T_40; // @[ALU.scala 38:20:@35.4]
	  wire  _T_42; // @[ALU.scala 39:20:@36.4]
	  wire  _T_44; // @[ALU.scala 40:20:@37.4]
	  wire  _T_46; // @[ALU.scala 41:20:@38.4]
	  wire  _T_48; // @[ALU.scala 42:20:@39.4]
	  wire [63:0] _T_49; // @[Mux.scala 61:16:@40.4]
	  wire [63:0] _T_50; // @[Mux.scala 61:16:@41.4]
	  wire [63:0] _T_51; // @[Mux.scala 61:16:@42.4]
	  wire [63:0] _T_52; // @[Mux.scala 61:16:@43.4]
	  wire [63:0] _T_53; // @[Mux.scala 61:16:@44.4]
	  wire [63:0] _T_54; // @[Mux.scala 61:16:@45.4]
	  wire [63:0] _T_55; // @[Mux.scala 61:16:@46.4]
	  wire [63:0] _T_56; // @[Mux.scala 61:16:@47.4]
	  assign _T_15 = io_opcode[4]; // @[ALUop.scala 20:29:@8.4]
	  assign _T_16 = ~ io_in2; // @[ALU.scala 19:54:@9.4]
	  assign _T_18 = _T_16 + 64'h1; // @[ALU.scala 19:62:@10.4]
	  assign _T_19 = _T_18[63:0]; // @[ALU.scala 19:62:@11.4]
	  assign _T_20 = _T_15 ? _T_19 : io_in2; // @[ALU.scala 19:35:@12.4]
	  assign add_result = io_in1 + _T_20; // @[ALU.scala 19:29:@13.4]
	  assign xor_result = io_in1 ^ io_in2; // @[ALU.scala 20:29:@14.4]
	  assign or_result = io_in1 | io_in2; // @[ALU.scala 21:29:@15.4]
	  assign and_result = io_in1 & io_in2; // @[ALU.scala 22:29:@16.4]
	  assign _T_21 = add_result[64]; // @[ALU.scala 24:41:@17.4]
	  assign sltu_result = ~ _T_21; // @[ALU.scala 24:30:@18.4]
	  assign _T_22 = xor_result[63]; // @[ALU.scala 25:40:@19.4]
	  assign slt_result = _T_22 ^ sltu_result; // @[ALU.scala 25:51:@20.4]
	  assign shamt = io_in2[4:0]; // @[ALU.scala 28:23:@21.4]
	  assign _GEN_0 = {{31'd0}, io_in1}; // @[ALU.scala 29:30:@22.4]
	  assign _T_23 = _GEN_0 << shamt; // @[ALU.scala 29:30:@22.4]
	  assign sll_result = _T_23[63:0]; // @[ALU.scala 29:39:@23.4]
	  assign _T_24 = $signed(io_in1); // @[ALU.scala 30:36:@24.4]
	  assign _T_25 = $signed(_T_24) >>> shamt; // @[ALU.scala 30:39:@25.4]
	  assign sra_result = $unsigned(_T_25); // @[ALU.scala 30:55:@26.4]
	  assign srl_result = io_in1 >> shamt; // @[ALU.scala 31:29:@27.4]
	  assign _T_26 = add_result[63:0]; // @[ALU.scala 33:33:@28.4]
	  assign _T_28 = io_opcode == 6'h12; // @[ALU.scala 34:20:@29.4]
	  assign _T_30 = {63'h0,sltu_result}; // @[Cat.scala 30:58:@30.4]
	  assign _T_32 = io_opcode == 6'h11; // @[ALU.scala 35:20:@31.4]
	  assign _T_34 = {63'h0,slt_result}; // @[Cat.scala 30:58:@32.4]
	  assign _T_36 = io_opcode == 6'h1; // @[ALU.scala 36:20:@33.4]
	  assign _T_38 = io_opcode == 6'h2; // @[ALU.scala 37:20:@34.4]
	  assign _T_40 = io_opcode == 6'h3; // @[ALU.scala 38:20:@35.4]
	  assign _T_42 = io_opcode == 6'h4; // @[ALU.scala 39:20:@36.4]
	  assign _T_44 = io_opcode == 6'h6; // @[ALU.scala 40:20:@37.4]
	  assign _T_46 = io_opcode == 6'h5; // @[ALU.scala 41:20:@38.4]
	  assign _T_48 = io_opcode == 6'h8; // @[ALU.scala 42:20:@39.4]
	  assign _T_49 = _T_48 ? io_in1 : _T_26; // @[Mux.scala 61:16:@40.4]
	  assign _T_50 = _T_46 ? srl_result : _T_49; // @[Mux.scala 61:16:@41.4]
	  assign _T_51 = _T_44 ? sra_result : _T_50; // @[Mux.scala 61:16:@42.4]
	  assign _T_52 = _T_42 ? sll_result : _T_51; // @[Mux.scala 61:16:@43.4]
	  assign _T_53 = _T_40 ? and_result : _T_52; // @[Mux.scala 61:16:@44.4]
	  assign _T_54 = _T_38 ? or_result : _T_53; // @[Mux.scala 61:16:@45.4]
	  assign _T_55 = _T_36 ? xor_result : _T_54; // @[Mux.scala 61:16:@46.4]
	  assign _T_56 = _T_32 ? _T_34 : _T_55; // @[Mux.scala 61:16:@47.4]
	  assign io_out = _T_28 ? _T_30 : _T_56; // @[ALU.scala 33:12:@49.4]
	  assign io_zero = io_out == 64'h0; // @[ALU.scala 45:13:@52.4]
	endmodule
	module IDU( // @[:@54.2]
%000042	  input  [31:0] io_inst, // @[:@57.4]
%000003	  output [3:0]  io_br_type, // @[:@57.4]
%000000	  output [1:0]  io_op1_sel, // @[:@57.4]
%000002	  output [1:0]  io_op2_sel, // @[:@57.4]
%000002	  output [5:0]  io_alu_op, // @[:@57.4]
%000001	  output [1:0]  io_wb_sel, // @[:@57.4]
%000001	  output        io_rf_wen, // @[:@57.4]
%000000	  output        io_mem_en, // @[:@57.4]
%000000	  output        io_mem_fcn, // @[:@57.4]
%000000	  output [2:0]  io_mem_msk // @[:@57.4]
	);
	  wire [31:0] _T_88; // @[Lookup.scala 9:38:@59.4]
	  wire  _T_89; // @[Lookup.scala 9:38:@60.4]
	  wire  _T_93; // @[Lookup.scala 9:38:@62.4]
	  wire  _T_97; // @[Lookup.scala 9:38:@64.4]
	  wire  _T_101; // @[Lookup.scala 9:38:@66.4]
	  wire  _T_105; // @[Lookup.scala 9:38:@68.4]
	  wire  _T_109; // @[Lookup.scala 9:38:@70.4]
	  wire  _T_113; // @[Lookup.scala 9:38:@72.4]
	  wire [31:0] _T_116; // @[Lookup.scala 9:38:@73.4]
	  wire  _T_117; // @[Lookup.scala 9:38:@74.4]
	  wire  _T_121; // @[Lookup.scala 9:38:@76.4]
	  wire  _T_125; // @[Lookup.scala 9:38:@78.4]
	  wire  _T_129; // @[Lookup.scala 9:38:@80.4]
	  wire  _T_133; // @[Lookup.scala 9:38:@82.4]
	  wire  _T_137; // @[Lookup.scala 9:38:@84.4]
	  wire  _T_141; // @[Lookup.scala 9:38:@86.4]
	  wire  _T_145; // @[Lookup.scala 9:38:@88.4]
	  wire [31:0] _T_148; // @[Lookup.scala 9:38:@89.4]
	  wire  _T_149; // @[Lookup.scala 9:38:@90.4]
	  wire  _T_153; // @[Lookup.scala 9:38:@92.4]
	  wire  _T_157; // @[Lookup.scala 9:38:@94.4]
	  wire [31:0] _T_160; // @[Lookup.scala 9:38:@95.4]
	  wire  _T_161; // @[Lookup.scala 9:38:@96.4]
	  wire  _T_165; // @[Lookup.scala 9:38:@98.4]
	  wire  _T_169; // @[Lookup.scala 9:38:@100.4]
	  wire  _T_173; // @[Lookup.scala 9:38:@102.4]
	  wire  _T_177; // @[Lookup.scala 9:38:@104.4]
	  wire  _T_181; // @[Lookup.scala 9:38:@106.4]
	  wire  _T_185; // @[Lookup.scala 9:38:@108.4]
	  wire  _T_189; // @[Lookup.scala 9:38:@110.4]
	  wire  _T_193; // @[Lookup.scala 9:38:@112.4]
	  wire  _T_197; // @[Lookup.scala 9:38:@114.4]
	  wire  _T_201; // @[Lookup.scala 9:38:@116.4]
	  wire  _T_205; // @[Lookup.scala 9:38:@118.4]
	  wire  _T_209; // @[Lookup.scala 9:38:@120.4]
	  wire  _T_213; // @[Lookup.scala 9:38:@122.4]
	  wire  _T_217; // @[Lookup.scala 9:38:@124.4]
	  wire  _T_221; // @[Lookup.scala 9:38:@126.4]
	  wire  _T_225; // @[Lookup.scala 9:38:@128.4]
	  wire  _T_229; // @[Lookup.scala 9:38:@130.4]
	  wire  _T_233; // @[Lookup.scala 9:38:@132.4]
	  wire  _T_237; // @[Lookup.scala 9:38:@134.4]
	  wire  _T_241; // @[Lookup.scala 9:38:@136.4]
	  wire  _T_245; // @[Lookup.scala 9:38:@138.4]
	  wire  _T_249; // @[Lookup.scala 9:38:@140.4]
	  wire  _T_253; // @[Lookup.scala 9:38:@142.4]
	  wire  _T_257; // @[Lookup.scala 9:38:@144.4]
	  wire  _T_261; // @[Lookup.scala 9:38:@146.4]
	  wire  _T_265; // @[Lookup.scala 9:38:@148.4]
	  wire  _T_269; // @[Lookup.scala 9:38:@150.4]
	  wire  _T_273; // @[Lookup.scala 9:38:@152.4]
	  wire  _T_277; // @[Lookup.scala 9:38:@154.4]
	  wire  _T_281; // @[Lookup.scala 9:38:@156.4]
	  wire [3:0] _T_343; // @[Lookup.scala 11:37:@219.4]
	  wire [3:0] _T_344; // @[Lookup.scala 11:37:@220.4]
	  wire [3:0] _T_345; // @[Lookup.scala 11:37:@221.4]
	  wire [3:0] _T_346; // @[Lookup.scala 11:37:@222.4]
	  wire [3:0] _T_347; // @[Lookup.scala 11:37:@223.4]
	  wire [3:0] _T_348; // @[Lookup.scala 11:37:@224.4]
	  wire [3:0] _T_349; // @[Lookup.scala 11:37:@225.4]
	  wire [3:0] _T_350; // @[Lookup.scala 11:37:@226.4]
	  wire [3:0] _T_351; // @[Lookup.scala 11:37:@227.4]
	  wire [3:0] _T_352; // @[Lookup.scala 11:37:@228.4]
	  wire [3:0] _T_353; // @[Lookup.scala 11:37:@229.4]
	  wire [3:0] _T_354; // @[Lookup.scala 11:37:@230.4]
	  wire [3:0] _T_355; // @[Lookup.scala 11:37:@231.4]
	  wire [3:0] _T_356; // @[Lookup.scala 11:37:@232.4]
	  wire [3:0] _T_357; // @[Lookup.scala 11:37:@233.4]
	  wire [3:0] _T_358; // @[Lookup.scala 11:37:@234.4]
	  wire [3:0] _T_359; // @[Lookup.scala 11:37:@235.4]
	  wire [3:0] _T_360; // @[Lookup.scala 11:37:@236.4]
	  wire [3:0] _T_361; // @[Lookup.scala 11:37:@237.4]
	  wire [3:0] _T_362; // @[Lookup.scala 11:37:@238.4]
	  wire [3:0] _T_363; // @[Lookup.scala 11:37:@239.4]
	  wire [3:0] _T_364; // @[Lookup.scala 11:37:@240.4]
	  wire [3:0] _T_365; // @[Lookup.scala 11:37:@241.4]
	  wire [3:0] _T_366; // @[Lookup.scala 11:37:@242.4]
	  wire [3:0] _T_367; // @[Lookup.scala 11:37:@243.4]
	  wire [3:0] _T_368; // @[Lookup.scala 11:37:@244.4]
	  wire [3:0] _T_369; // @[Lookup.scala 11:37:@245.4]
	  wire [3:0] _T_370; // @[Lookup.scala 11:37:@246.4]
	  wire [3:0] _T_371; // @[Lookup.scala 11:37:@247.4]
	  wire [3:0] _T_372; // @[Lookup.scala 11:37:@248.4]
	  wire [3:0] _T_373; // @[Lookup.scala 11:37:@249.4]
	  wire [3:0] _T_374; // @[Lookup.scala 11:37:@250.4]
	  wire [3:0] _T_375; // @[Lookup.scala 11:37:@251.4]
	  wire [3:0] _T_376; // @[Lookup.scala 11:37:@252.4]
	  wire [3:0] _T_377; // @[Lookup.scala 11:37:@253.4]
	  wire [1:0] _T_388; // @[Lookup.scala 11:37:@265.4]
	  wire [1:0] _T_389; // @[Lookup.scala 11:37:@266.4]
	  wire [1:0] _T_390; // @[Lookup.scala 11:37:@267.4]
	  wire [1:0] _T_391; // @[Lookup.scala 11:37:@268.4]
	  wire [1:0] _T_392; // @[Lookup.scala 11:37:@269.4]
	  wire [1:0] _T_393; // @[Lookup.scala 11:37:@270.4]
	  wire [1:0] _T_394; // @[Lookup.scala 11:37:@271.4]
	  wire [1:0] _T_395; // @[Lookup.scala 11:37:@272.4]
	  wire [1:0] _T_396; // @[Lookup.scala 11:37:@273.4]
	  wire [1:0] _T_397; // @[Lookup.scala 11:37:@274.4]
	  wire [1:0] _T_398; // @[Lookup.scala 11:37:@275.4]
	  wire [1:0] _T_399; // @[Lookup.scala 11:37:@276.4]
	  wire [1:0] _T_400; // @[Lookup.scala 11:37:@277.4]
	  wire [1:0] _T_401; // @[Lookup.scala 11:37:@278.4]
	  wire [1:0] _T_402; // @[Lookup.scala 11:37:@279.4]
	  wire [1:0] _T_403; // @[Lookup.scala 11:37:@280.4]
	  wire [1:0] _T_404; // @[Lookup.scala 11:37:@281.4]
	  wire [1:0] _T_405; // @[Lookup.scala 11:37:@282.4]
	  wire [1:0] _T_406; // @[Lookup.scala 11:37:@283.4]
	  wire [1:0] _T_407; // @[Lookup.scala 11:37:@284.4]
	  wire [1:0] _T_408; // @[Lookup.scala 11:37:@285.4]
	  wire [1:0] _T_409; // @[Lookup.scala 11:37:@286.4]
	  wire [1:0] _T_410; // @[Lookup.scala 11:37:@287.4]
	  wire [1:0] _T_411; // @[Lookup.scala 11:37:@288.4]
	  wire [1:0] _T_412; // @[Lookup.scala 11:37:@289.4]
	  wire [1:0] _T_413; // @[Lookup.scala 11:37:@290.4]
	  wire [1:0] _T_414; // @[Lookup.scala 11:37:@291.4]
	  wire [1:0] _T_415; // @[Lookup.scala 11:37:@292.4]
	  wire [1:0] _T_416; // @[Lookup.scala 11:37:@293.4]
	  wire [1:0] _T_417; // @[Lookup.scala 11:37:@294.4]
	  wire [1:0] _T_418; // @[Lookup.scala 11:37:@295.4]
	  wire [1:0] _T_419; // @[Lookup.scala 11:37:@296.4]
	  wire [1:0] _T_420; // @[Lookup.scala 11:37:@297.4]
	  wire [1:0] _T_421; // @[Lookup.scala 11:37:@298.4]
	  wire [1:0] _T_422; // @[Lookup.scala 11:37:@299.4]
	  wire [1:0] _T_423; // @[Lookup.scala 11:37:@300.4]
	  wire [1:0] _T_424; // @[Lookup.scala 11:37:@301.4]
	  wire [1:0] _T_425; // @[Lookup.scala 11:37:@302.4]
	  wire [1:0] _T_445; // @[Lookup.scala 11:37:@323.4]
	  wire [1:0] _T_446; // @[Lookup.scala 11:37:@324.4]
	  wire [1:0] _T_447; // @[Lookup.scala 11:37:@325.4]
	  wire [1:0] _T_448; // @[Lookup.scala 11:37:@326.4]
	  wire [1:0] _T_449; // @[Lookup.scala 11:37:@327.4]
	  wire [1:0] _T_450; // @[Lookup.scala 11:37:@328.4]
	  wire [1:0] _T_451; // @[Lookup.scala 11:37:@329.4]
	  wire [1:0] _T_452; // @[Lookup.scala 11:37:@330.4]
	  wire [1:0] _T_453; // @[Lookup.scala 11:37:@331.4]
	  wire [1:0] _T_454; // @[Lookup.scala 11:37:@332.4]
	  wire [1:0] _T_455; // @[Lookup.scala 11:37:@333.4]
	  wire [1:0] _T_456; // @[Lookup.scala 11:37:@334.4]
	  wire [1:0] _T_457; // @[Lookup.scala 11:37:@335.4]
	  wire [1:0] _T_458; // @[Lookup.scala 11:37:@336.4]
	  wire [1:0] _T_459; // @[Lookup.scala 11:37:@337.4]
	  wire [1:0] _T_460; // @[Lookup.scala 11:37:@338.4]
	  wire [1:0] _T_461; // @[Lookup.scala 11:37:@339.4]
	  wire [1:0] _T_462; // @[Lookup.scala 11:37:@340.4]
	  wire [1:0] _T_463; // @[Lookup.scala 11:37:@341.4]
	  wire [1:0] _T_464; // @[Lookup.scala 11:37:@342.4]
	  wire [1:0] _T_465; // @[Lookup.scala 11:37:@343.4]
	  wire [1:0] _T_466; // @[Lookup.scala 11:37:@344.4]
	  wire [1:0] _T_467; // @[Lookup.scala 11:37:@345.4]
	  wire [1:0] _T_468; // @[Lookup.scala 11:37:@346.4]
	  wire [1:0] _T_469; // @[Lookup.scala 11:37:@347.4]
	  wire [1:0] _T_470; // @[Lookup.scala 11:37:@348.4]
	  wire [1:0] _T_471; // @[Lookup.scala 11:37:@349.4]
	  wire [1:0] _T_472; // @[Lookup.scala 11:37:@350.4]
	  wire [1:0] _T_473; // @[Lookup.scala 11:37:@351.4]
	  wire [3:0] _T_481; // @[Lookup.scala 11:37:@360.4]
	  wire [3:0] _T_482; // @[Lookup.scala 11:37:@361.4]
	  wire [3:0] _T_483; // @[Lookup.scala 11:37:@362.4]
	  wire [3:0] _T_484; // @[Lookup.scala 11:37:@363.4]
	  wire [3:0] _T_485; // @[Lookup.scala 11:37:@364.4]
	  wire [3:0] _T_486; // @[Lookup.scala 11:37:@365.4]
	  wire [4:0] _T_487; // @[Lookup.scala 11:37:@366.4]
	  wire [4:0] _T_488; // @[Lookup.scala 11:37:@367.4]
	  wire [4:0] _T_489; // @[Lookup.scala 11:37:@368.4]
	  wire [4:0] _T_490; // @[Lookup.scala 11:37:@369.4]
	  wire [4:0] _T_491; // @[Lookup.scala 11:37:@370.4]
	  wire [4:0] _T_492; // @[Lookup.scala 11:37:@371.4]
	  wire [4:0] _T_493; // @[Lookup.scala 11:37:@372.4]
	  wire [4:0] _T_494; // @[Lookup.scala 11:37:@373.4]
	  wire [4:0] _T_495; // @[Lookup.scala 11:37:@374.4]
	  wire [4:0] _T_496; // @[Lookup.scala 11:37:@375.4]
	  wire [4:0] _T_497; // @[Lookup.scala 11:37:@376.4]
	  wire [4:0] _T_498; // @[Lookup.scala 11:37:@377.4]
	  wire [4:0] _T_499; // @[Lookup.scala 11:37:@378.4]
	  wire [4:0] _T_500; // @[Lookup.scala 11:37:@379.4]
	  wire [4:0] _T_501; // @[Lookup.scala 11:37:@380.4]
	  wire [4:0] _T_502; // @[Lookup.scala 11:37:@381.4]
	  wire [4:0] _T_503; // @[Lookup.scala 11:37:@382.4]
	  wire [4:0] _T_504; // @[Lookup.scala 11:37:@383.4]
	  wire [4:0] _T_505; // @[Lookup.scala 11:37:@384.4]
	  wire [4:0] _T_506; // @[Lookup.scala 11:37:@385.4]
	  wire [4:0] _T_507; // @[Lookup.scala 11:37:@386.4]
	  wire [4:0] _T_508; // @[Lookup.scala 11:37:@387.4]
	  wire [4:0] _T_509; // @[Lookup.scala 11:37:@388.4]
	  wire [4:0] _T_510; // @[Lookup.scala 11:37:@389.4]
	  wire [4:0] _T_511; // @[Lookup.scala 11:37:@390.4]
	  wire [4:0] _T_512; // @[Lookup.scala 11:37:@391.4]
	  wire [4:0] _T_513; // @[Lookup.scala 11:37:@392.4]
	  wire [4:0] _T_514; // @[Lookup.scala 11:37:@393.4]
	  wire [4:0] _T_515; // @[Lookup.scala 11:37:@394.4]
	  wire [4:0] _T_516; // @[Lookup.scala 11:37:@395.4]
	  wire [4:0] _T_517; // @[Lookup.scala 11:37:@396.4]
	  wire [4:0] _T_518; // @[Lookup.scala 11:37:@397.4]
	  wire [4:0] _T_519; // @[Lookup.scala 11:37:@398.4]
	  wire [4:0] _T_520; // @[Lookup.scala 11:37:@399.4]
	  wire [4:0] _T_521; // @[Lookup.scala 11:37:@400.4]
%000002	  wire [4:0] csignals_4; // @[Lookup.scala 11:37:@401.4]
	  wire [1:0] _T_529; // @[Lookup.scala 11:37:@409.4]
	  wire [1:0] _T_530; // @[Lookup.scala 11:37:@410.4]
	  wire [1:0] _T_531; // @[Lookup.scala 11:37:@411.4]
	  wire [1:0] _T_532; // @[Lookup.scala 11:37:@412.4]
	  wire [1:0] _T_533; // @[Lookup.scala 11:37:@413.4]
	  wire [1:0] _T_534; // @[Lookup.scala 11:37:@414.4]
	  wire [1:0] _T_535; // @[Lookup.scala 11:37:@415.4]
	  wire [1:0] _T_536; // @[Lookup.scala 11:37:@416.4]
	  wire [1:0] _T_537; // @[Lookup.scala 11:37:@417.4]
	  wire [1:0] _T_538; // @[Lookup.scala 11:37:@418.4]
	  wire [1:0] _T_539; // @[Lookup.scala 11:37:@419.4]
	  wire [1:0] _T_540; // @[Lookup.scala 11:37:@420.4]
	  wire [1:0] _T_541; // @[Lookup.scala 11:37:@421.4]
	  wire [1:0] _T_542; // @[Lookup.scala 11:37:@422.4]
	  wire [1:0] _T_543; // @[Lookup.scala 11:37:@423.4]
	  wire [1:0] _T_544; // @[Lookup.scala 11:37:@424.4]
	  wire [1:0] _T_545; // @[Lookup.scala 11:37:@425.4]
	  wire [1:0] _T_546; // @[Lookup.scala 11:37:@426.4]
	  wire [1:0] _T_547; // @[Lookup.scala 11:37:@427.4]
	  wire [1:0] _T_548; // @[Lookup.scala 11:37:@428.4]
	  wire [1:0] _T_549; // @[Lookup.scala 11:37:@429.4]
	  wire [1:0] _T_550; // @[Lookup.scala 11:37:@430.4]
	  wire [1:0] _T_551; // @[Lookup.scala 11:37:@431.4]
	  wire [1:0] _T_552; // @[Lookup.scala 11:37:@432.4]
	  wire [1:0] _T_553; // @[Lookup.scala 11:37:@433.4]
	  wire [1:0] _T_554; // @[Lookup.scala 11:37:@434.4]
	  wire [1:0] _T_555; // @[Lookup.scala 11:37:@435.4]
	  wire [1:0] _T_556; // @[Lookup.scala 11:37:@436.4]
	  wire [1:0] _T_557; // @[Lookup.scala 11:37:@437.4]
	  wire [1:0] _T_558; // @[Lookup.scala 11:37:@438.4]
	  wire [1:0] _T_559; // @[Lookup.scala 11:37:@439.4]
	  wire [1:0] _T_560; // @[Lookup.scala 11:37:@440.4]
	  wire [1:0] _T_561; // @[Lookup.scala 11:37:@441.4]
	  wire [1:0] _T_562; // @[Lookup.scala 11:37:@442.4]
	  wire [1:0] _T_563; // @[Lookup.scala 11:37:@443.4]
	  wire [1:0] _T_564; // @[Lookup.scala 11:37:@444.4]
	  wire [1:0] _T_565; // @[Lookup.scala 11:37:@445.4]
	  wire [1:0] _T_566; // @[Lookup.scala 11:37:@446.4]
	  wire [1:0] _T_567; // @[Lookup.scala 11:37:@447.4]
	  wire [1:0] _T_568; // @[Lookup.scala 11:37:@448.4]
	  wire [1:0] _T_569; // @[Lookup.scala 11:37:@449.4]
	  wire  _T_578; // @[Lookup.scala 11:37:@459.4]
	  wire  _T_579; // @[Lookup.scala 11:37:@460.4]
	  wire  _T_580; // @[Lookup.scala 11:37:@461.4]
	  wire  _T_581; // @[Lookup.scala 11:37:@462.4]
	  wire  _T_582; // @[Lookup.scala 11:37:@463.4]
	  wire  _T_583; // @[Lookup.scala 11:37:@464.4]
	  wire  _T_584; // @[Lookup.scala 11:37:@465.4]
	  wire  _T_585; // @[Lookup.scala 11:37:@466.4]
	  wire  _T_586; // @[Lookup.scala 11:37:@467.4]
	  wire  _T_587; // @[Lookup.scala 11:37:@468.4]
	  wire  _T_588; // @[Lookup.scala 11:37:@469.4]
	  wire  _T_589; // @[Lookup.scala 11:37:@470.4]
	  wire  _T_590; // @[Lookup.scala 11:37:@471.4]
	  wire  _T_591; // @[Lookup.scala 11:37:@472.4]
	  wire  _T_592; // @[Lookup.scala 11:37:@473.4]
	  wire  _T_593; // @[Lookup.scala 11:37:@474.4]
	  wire  _T_594; // @[Lookup.scala 11:37:@475.4]
	  wire  _T_595; // @[Lookup.scala 11:37:@476.4]
	  wire  _T_596; // @[Lookup.scala 11:37:@477.4]
	  wire  _T_597; // @[Lookup.scala 11:37:@478.4]
	  wire  _T_598; // @[Lookup.scala 11:37:@479.4]
	  wire  _T_599; // @[Lookup.scala 11:37:@480.4]
	  wire  _T_600; // @[Lookup.scala 11:37:@481.4]
	  wire  _T_601; // @[Lookup.scala 11:37:@482.4]
	  wire  _T_602; // @[Lookup.scala 11:37:@483.4]
	  wire  _T_603; // @[Lookup.scala 11:37:@484.4]
	  wire  _T_604; // @[Lookup.scala 11:37:@485.4]
	  wire  _T_605; // @[Lookup.scala 11:37:@486.4]
	  wire  _T_606; // @[Lookup.scala 11:37:@487.4]
	  wire  _T_607; // @[Lookup.scala 11:37:@488.4]
	  wire  _T_608; // @[Lookup.scala 11:37:@489.4]
	  wire  _T_609; // @[Lookup.scala 11:37:@490.4]
	  wire  _T_610; // @[Lookup.scala 11:37:@491.4]
	  wire  _T_611; // @[Lookup.scala 11:37:@492.4]
	  wire  _T_612; // @[Lookup.scala 11:37:@493.4]
	  wire  _T_613; // @[Lookup.scala 11:37:@494.4]
	  wire  _T_614; // @[Lookup.scala 11:37:@495.4]
	  wire  _T_615; // @[Lookup.scala 11:37:@496.4]
	  wire  _T_616; // @[Lookup.scala 11:37:@497.4]
	  wire  _T_617; // @[Lookup.scala 11:37:@498.4]
	  wire  _T_619; // @[Lookup.scala 11:37:@501.4]
	  wire  _T_620; // @[Lookup.scala 11:37:@502.4]
	  wire  _T_621; // @[Lookup.scala 11:37:@503.4]
	  wire  _T_622; // @[Lookup.scala 11:37:@504.4]
	  wire  _T_623; // @[Lookup.scala 11:37:@505.4]
	  wire  _T_624; // @[Lookup.scala 11:37:@506.4]
	  wire  _T_625; // @[Lookup.scala 11:37:@507.4]
	  wire  _T_626; // @[Lookup.scala 11:37:@508.4]
	  wire  _T_627; // @[Lookup.scala 11:37:@509.4]
	  wire  _T_628; // @[Lookup.scala 11:37:@510.4]
	  wire  _T_629; // @[Lookup.scala 11:37:@511.4]
	  wire  _T_630; // @[Lookup.scala 11:37:@512.4]
	  wire  _T_631; // @[Lookup.scala 11:37:@513.4]
	  wire  _T_632; // @[Lookup.scala 11:37:@514.4]
	  wire  _T_633; // @[Lookup.scala 11:37:@515.4]
	  wire  _T_634; // @[Lookup.scala 11:37:@516.4]
	  wire  _T_635; // @[Lookup.scala 11:37:@517.4]
	  wire  _T_636; // @[Lookup.scala 11:37:@518.4]
	  wire  _T_637; // @[Lookup.scala 11:37:@519.4]
	  wire  _T_638; // @[Lookup.scala 11:37:@520.4]
	  wire  _T_639; // @[Lookup.scala 11:37:@521.4]
	  wire  _T_640; // @[Lookup.scala 11:37:@522.4]
	  wire  _T_641; // @[Lookup.scala 11:37:@523.4]
	  wire  _T_642; // @[Lookup.scala 11:37:@524.4]
	  wire  _T_643; // @[Lookup.scala 11:37:@525.4]
	  wire  _T_644; // @[Lookup.scala 11:37:@526.4]
	  wire  _T_645; // @[Lookup.scala 11:37:@527.4]
	  wire  _T_646; // @[Lookup.scala 11:37:@528.4]
	  wire  _T_647; // @[Lookup.scala 11:37:@529.4]
	  wire  _T_648; // @[Lookup.scala 11:37:@530.4]
	  wire  _T_649; // @[Lookup.scala 11:37:@531.4]
	  wire  _T_650; // @[Lookup.scala 11:37:@532.4]
	  wire  _T_651; // @[Lookup.scala 11:37:@533.4]
	  wire  _T_652; // @[Lookup.scala 11:37:@534.4]
	  wire  _T_653; // @[Lookup.scala 11:37:@535.4]
	  wire  _T_654; // @[Lookup.scala 11:37:@536.4]
	  wire  _T_655; // @[Lookup.scala 11:37:@537.4]
	  wire  _T_656; // @[Lookup.scala 11:37:@538.4]
	  wire  _T_657; // @[Lookup.scala 11:37:@539.4]
	  wire  _T_658; // @[Lookup.scala 11:37:@540.4]
	  wire  _T_659; // @[Lookup.scala 11:37:@541.4]
	  wire  _T_660; // @[Lookup.scala 11:37:@542.4]
	  wire  _T_661; // @[Lookup.scala 11:37:@543.4]
	  wire  _T_662; // @[Lookup.scala 11:37:@544.4]
	  wire  _T_663; // @[Lookup.scala 11:37:@545.4]
	  wire  _T_664; // @[Lookup.scala 11:37:@546.4]
	  wire  _T_665; // @[Lookup.scala 11:37:@547.4]
	  wire  _T_709; // @[Lookup.scala 11:37:@592.4]
	  wire  _T_710; // @[Lookup.scala 11:37:@593.4]
	  wire  _T_711; // @[Lookup.scala 11:37:@594.4]
	  wire  _T_712; // @[Lookup.scala 11:37:@595.4]
	  wire  _T_713; // @[Lookup.scala 11:37:@596.4]
	  wire [2:0] _T_756; // @[Lookup.scala 11:37:@640.4]
	  wire [2:0] _T_757; // @[Lookup.scala 11:37:@641.4]
	  wire [2:0] _T_758; // @[Lookup.scala 11:37:@642.4]
	  wire [2:0] _T_759; // @[Lookup.scala 11:37:@643.4]
	  wire [2:0] _T_760; // @[Lookup.scala 11:37:@644.4]
	  wire [2:0] _T_761; // @[Lookup.scala 11:37:@645.4]
	  assign _T_88 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@59.4]
	  assign _T_89 = 32'h2003 == _T_88; // @[Lookup.scala 9:38:@60.4]
	  assign _T_93 = 32'h3 == _T_88; // @[Lookup.scala 9:38:@62.4]
	  assign _T_97 = 32'h4003 == _T_88; // @[Lookup.scala 9:38:@64.4]
	  assign _T_101 = 32'h5003 == _T_88; // @[Lookup.scala 9:38:@66.4]
	  assign _T_105 = 32'h2023 == _T_88; // @[Lookup.scala 9:38:@68.4]
	  assign _T_109 = 32'h23 == _T_88; // @[Lookup.scala 9:38:@70.4]
	  assign _T_113 = 32'h1023 == _T_88; // @[Lookup.scala 9:38:@72.4]
	  assign _T_116 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@73.4]
	  assign _T_117 = 32'h17 == _T_116; // @[Lookup.scala 9:38:@74.4]
	  assign _T_121 = 32'h37 == _T_116; // @[Lookup.scala 9:38:@76.4]
	  assign _T_125 = 32'h13 == _T_88; // @[Lookup.scala 9:38:@78.4]
	  assign _T_129 = 32'h7013 == _T_88; // @[Lookup.scala 9:38:@80.4]
	  assign _T_133 = 32'h6013 == _T_88; // @[Lookup.scala 9:38:@82.4]
	  assign _T_137 = 32'h4013 == _T_88; // @[Lookup.scala 9:38:@84.4]
	  assign _T_141 = 32'h2013 == _T_88; // @[Lookup.scala 9:38:@86.4]
	  assign _T_145 = 32'h3013 == _T_88; // @[Lookup.scala 9:38:@88.4]
	  assign _T_148 = io_inst & 32'hfc00707f; // @[Lookup.scala 9:38:@89.4]
	  assign _T_149 = 32'h1013 == _T_148; // @[Lookup.scala 9:38:@90.4]
	  assign _T_153 = 32'h40005013 == _T_148; // @[Lookup.scala 9:38:@92.4]
	  assign _T_157 = 32'h5013 == _T_148; // @[Lookup.scala 9:38:@94.4]
	  assign _T_160 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@95.4]
	  assign _T_161 = 32'h1033 == _T_160; // @[Lookup.scala 9:38:@96.4]
	  assign _T_165 = 32'h33 == _T_160; // @[Lookup.scala 9:38:@98.4]
	  assign _T_169 = 32'h40000033 == _T_160; // @[Lookup.scala 9:38:@100.4]
	  assign _T_173 = 32'h2033 == _T_160; // @[Lookup.scala 9:38:@102.4]
	  assign _T_177 = 32'h3033 == _T_160; // @[Lookup.scala 9:38:@104.4]
	  assign _T_181 = 32'h7033 == _T_160; // @[Lookup.scala 9:38:@106.4]
	  assign _T_185 = 32'h6033 == _T_160; // @[Lookup.scala 9:38:@108.4]
	  assign _T_189 = 32'h4033 == _T_160; // @[Lookup.scala 9:38:@110.4]
	  assign _T_193 = 32'h40005033 == _T_160; // @[Lookup.scala 9:38:@112.4]
	  assign _T_197 = 32'h5033 == _T_160; // @[Lookup.scala 9:38:@114.4]
	  assign _T_201 = 32'h6f == _T_116; // @[Lookup.scala 9:38:@116.4]
	  assign _T_205 = 32'h67 == _T_88; // @[Lookup.scala 9:38:@118.4]
	  assign _T_209 = 32'h63 == _T_88; // @[Lookup.scala 9:38:@120.4]
	  assign _T_213 = 32'h1063 == _T_88; // @[Lookup.scala 9:38:@122.4]
	  assign _T_217 = 32'h5063 == _T_88; // @[Lookup.scala 9:38:@124.4]
	  assign _T_221 = 32'h7063 == _T_88; // @[Lookup.scala 9:38:@126.4]
	  assign _T_225 = 32'h4063 == _T_88; // @[Lookup.scala 9:38:@128.4]
	  assign _T_229 = 32'h6063 == _T_88; // @[Lookup.scala 9:38:@130.4]
	  assign _T_233 = 32'h5073 == _T_88; // @[Lookup.scala 9:38:@132.4]
	  assign _T_237 = 32'h6073 == _T_88; // @[Lookup.scala 9:38:@134.4]
	  assign _T_241 = 32'h7073 == _T_88; // @[Lookup.scala 9:38:@136.4]
	  assign _T_245 = 32'h1073 == _T_88; // @[Lookup.scala 9:38:@138.4]
	  assign _T_249 = 32'h2073 == _T_88; // @[Lookup.scala 9:38:@140.4]
	  assign _T_253 = 32'h3073 == _T_88; // @[Lookup.scala 9:38:@142.4]
	  assign _T_257 = 32'h73 == io_inst; // @[Lookup.scala 9:38:@144.4]
	  assign _T_261 = 32'h30200073 == io_inst; // @[Lookup.scala 9:38:@146.4]
	  assign _T_265 = 32'h7b200073 == io_inst; // @[Lookup.scala 9:38:@148.4]
	  assign _T_269 = 32'h100073 == io_inst; // @[Lookup.scala 9:38:@150.4]
	  assign _T_273 = 32'h10500073 == io_inst; // @[Lookup.scala 9:38:@152.4]
	  assign _T_277 = 32'h100f == _T_88; // @[Lookup.scala 9:38:@154.4]
	  assign _T_281 = 32'hf == _T_88; // @[Lookup.scala 9:38:@156.4]
	  assign _T_343 = _T_229 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37:@219.4]
	  assign _T_344 = _T_225 ? 4'h5 : _T_343; // @[Lookup.scala 11:37:@220.4]
	  assign _T_345 = _T_221 ? 4'h4 : _T_344; // @[Lookup.scala 11:37:@221.4]
	  assign _T_346 = _T_217 ? 4'h3 : _T_345; // @[Lookup.scala 11:37:@222.4]
	  assign _T_347 = _T_213 ? 4'h1 : _T_346; // @[Lookup.scala 11:37:@223.4]
	  assign _T_348 = _T_209 ? 4'h2 : _T_347; // @[Lookup.scala 11:37:@224.4]
	  assign _T_349 = _T_205 ? 4'h8 : _T_348; // @[Lookup.scala 11:37:@225.4]
	  assign _T_350 = _T_201 ? 4'h7 : _T_349; // @[Lookup.scala 11:37:@226.4]
	  assign _T_351 = _T_197 ? 4'h0 : _T_350; // @[Lookup.scala 11:37:@227.4]
	  assign _T_352 = _T_193 ? 4'h0 : _T_351; // @[Lookup.scala 11:37:@228.4]
	  assign _T_353 = _T_189 ? 4'h0 : _T_352; // @[Lookup.scala 11:37:@229.4]
	  assign _T_354 = _T_185 ? 4'h0 : _T_353; // @[Lookup.scala 11:37:@230.4]
	  assign _T_355 = _T_181 ? 4'h0 : _T_354; // @[Lookup.scala 11:37:@231.4]
	  assign _T_356 = _T_177 ? 4'h0 : _T_355; // @[Lookup.scala 11:37:@232.4]
	  assign _T_357 = _T_173 ? 4'h0 : _T_356; // @[Lookup.scala 11:37:@233.4]
	  assign _T_358 = _T_169 ? 4'h0 : _T_357; // @[Lookup.scala 11:37:@234.4]
	  assign _T_359 = _T_165 ? 4'h0 : _T_358; // @[Lookup.scala 11:37:@235.4]
	  assign _T_360 = _T_161 ? 4'h0 : _T_359; // @[Lookup.scala 11:37:@236.4]
	  assign _T_361 = _T_157 ? 4'h0 : _T_360; // @[Lookup.scala 11:37:@237.4]
	  assign _T_362 = _T_153 ? 4'h0 : _T_361; // @[Lookup.scala 11:37:@238.4]
	  assign _T_363 = _T_149 ? 4'h0 : _T_362; // @[Lookup.scala 11:37:@239.4]
	  assign _T_364 = _T_145 ? 4'h0 : _T_363; // @[Lookup.scala 11:37:@240.4]
	  assign _T_365 = _T_141 ? 4'h0 : _T_364; // @[Lookup.scala 11:37:@241.4]
	  assign _T_366 = _T_137 ? 4'h0 : _T_365; // @[Lookup.scala 11:37:@242.4]
	  assign _T_367 = _T_133 ? 4'h0 : _T_366; // @[Lookup.scala 11:37:@243.4]
	  assign _T_368 = _T_129 ? 4'h0 : _T_367; // @[Lookup.scala 11:37:@244.4]
	  assign _T_369 = _T_125 ? 4'h0 : _T_368; // @[Lookup.scala 11:37:@245.4]
	  assign _T_370 = _T_121 ? 4'h0 : _T_369; // @[Lookup.scala 11:37:@246.4]
	  assign _T_371 = _T_117 ? 4'h0 : _T_370; // @[Lookup.scala 11:37:@247.4]
	  assign _T_372 = _T_113 ? 4'h0 : _T_371; // @[Lookup.scala 11:37:@248.4]
	  assign _T_373 = _T_109 ? 4'h0 : _T_372; // @[Lookup.scala 11:37:@249.4]
	  assign _T_374 = _T_105 ? 4'h0 : _T_373; // @[Lookup.scala 11:37:@250.4]
	  assign _T_375 = _T_101 ? 4'h0 : _T_374; // @[Lookup.scala 11:37:@251.4]
	  assign _T_376 = _T_97 ? 4'h0 : _T_375; // @[Lookup.scala 11:37:@252.4]
	  assign _T_377 = _T_93 ? 4'h0 : _T_376; // @[Lookup.scala 11:37:@253.4]
	  assign _T_388 = _T_241 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@265.4]
	  assign _T_389 = _T_237 ? 2'h2 : _T_388; // @[Lookup.scala 11:37:@266.4]
	  assign _T_390 = _T_233 ? 2'h2 : _T_389; // @[Lookup.scala 11:37:@267.4]
	  assign _T_391 = _T_229 ? 2'h0 : _T_390; // @[Lookup.scala 11:37:@268.4]
	  assign _T_392 = _T_225 ? 2'h0 : _T_391; // @[Lookup.scala 11:37:@269.4]
	  assign _T_393 = _T_221 ? 2'h0 : _T_392; // @[Lookup.scala 11:37:@270.4]
	  assign _T_394 = _T_217 ? 2'h0 : _T_393; // @[Lookup.scala 11:37:@271.4]
	  assign _T_395 = _T_213 ? 2'h0 : _T_394; // @[Lookup.scala 11:37:@272.4]
	  assign _T_396 = _T_209 ? 2'h0 : _T_395; // @[Lookup.scala 11:37:@273.4]
	  assign _T_397 = _T_205 ? 2'h0 : _T_396; // @[Lookup.scala 11:37:@274.4]
	  assign _T_398 = _T_201 ? 2'h0 : _T_397; // @[Lookup.scala 11:37:@275.4]
	  assign _T_399 = _T_197 ? 2'h0 : _T_398; // @[Lookup.scala 11:37:@276.4]
	  assign _T_400 = _T_193 ? 2'h0 : _T_399; // @[Lookup.scala 11:37:@277.4]
	  assign _T_401 = _T_189 ? 2'h0 : _T_400; // @[Lookup.scala 11:37:@278.4]
	  assign _T_402 = _T_185 ? 2'h0 : _T_401; // @[Lookup.scala 11:37:@279.4]
	  assign _T_403 = _T_181 ? 2'h0 : _T_402; // @[Lookup.scala 11:37:@280.4]
	  assign _T_404 = _T_177 ? 2'h0 : _T_403; // @[Lookup.scala 11:37:@281.4]
	  assign _T_405 = _T_173 ? 2'h0 : _T_404; // @[Lookup.scala 11:37:@282.4]
	  assign _T_406 = _T_169 ? 2'h0 : _T_405; // @[Lookup.scala 11:37:@283.4]
	  assign _T_407 = _T_165 ? 2'h0 : _T_406; // @[Lookup.scala 11:37:@284.4]
	  assign _T_408 = _T_161 ? 2'h0 : _T_407; // @[Lookup.scala 11:37:@285.4]
	  assign _T_409 = _T_157 ? 2'h0 : _T_408; // @[Lookup.scala 11:37:@286.4]
	  assign _T_410 = _T_153 ? 2'h0 : _T_409; // @[Lookup.scala 11:37:@287.4]
	  assign _T_411 = _T_149 ? 2'h0 : _T_410; // @[Lookup.scala 11:37:@288.4]
	  assign _T_412 = _T_145 ? 2'h0 : _T_411; // @[Lookup.scala 11:37:@289.4]
	  assign _T_413 = _T_141 ? 2'h0 : _T_412; // @[Lookup.scala 11:37:@290.4]
	  assign _T_414 = _T_137 ? 2'h0 : _T_413; // @[Lookup.scala 11:37:@291.4]
	  assign _T_415 = _T_133 ? 2'h0 : _T_414; // @[Lookup.scala 11:37:@292.4]
	  assign _T_416 = _T_129 ? 2'h0 : _T_415; // @[Lookup.scala 11:37:@293.4]
	  assign _T_417 = _T_125 ? 2'h0 : _T_416; // @[Lookup.scala 11:37:@294.4]
	  assign _T_418 = _T_121 ? 2'h1 : _T_417; // @[Lookup.scala 11:37:@295.4]
	  assign _T_419 = _T_117 ? 2'h1 : _T_418; // @[Lookup.scala 11:37:@296.4]
	  assign _T_420 = _T_113 ? 2'h0 : _T_419; // @[Lookup.scala 11:37:@297.4]
	  assign _T_421 = _T_109 ? 2'h0 : _T_420; // @[Lookup.scala 11:37:@298.4]
	  assign _T_422 = _T_105 ? 2'h0 : _T_421; // @[Lookup.scala 11:37:@299.4]
	  assign _T_423 = _T_101 ? 2'h0 : _T_422; // @[Lookup.scala 11:37:@300.4]
	  assign _T_424 = _T_97 ? 2'h0 : _T_423; // @[Lookup.scala 11:37:@301.4]
	  assign _T_425 = _T_93 ? 2'h0 : _T_424; // @[Lookup.scala 11:37:@302.4]
	  assign _T_445 = _T_205 ? 2'h1 : 2'h0; // @[Lookup.scala 11:37:@323.4]
	  assign _T_446 = _T_201 ? 2'h0 : _T_445; // @[Lookup.scala 11:37:@324.4]
	  assign _T_447 = _T_197 ? 2'h0 : _T_446; // @[Lookup.scala 11:37:@325.4]
	  assign _T_448 = _T_193 ? 2'h0 : _T_447; // @[Lookup.scala 11:37:@326.4]
	  assign _T_449 = _T_189 ? 2'h0 : _T_448; // @[Lookup.scala 11:37:@327.4]
	  assign _T_450 = _T_185 ? 2'h0 : _T_449; // @[Lookup.scala 11:37:@328.4]
	  assign _T_451 = _T_181 ? 2'h0 : _T_450; // @[Lookup.scala 11:37:@329.4]
	  assign _T_452 = _T_177 ? 2'h0 : _T_451; // @[Lookup.scala 11:37:@330.4]
	  assign _T_453 = _T_173 ? 2'h0 : _T_452; // @[Lookup.scala 11:37:@331.4]
	  assign _T_454 = _T_169 ? 2'h0 : _T_453; // @[Lookup.scala 11:37:@332.4]
	  assign _T_455 = _T_165 ? 2'h0 : _T_454; // @[Lookup.scala 11:37:@333.4]
	  assign _T_456 = _T_161 ? 2'h0 : _T_455; // @[Lookup.scala 11:37:@334.4]
	  assign _T_457 = _T_157 ? 2'h1 : _T_456; // @[Lookup.scala 11:37:@335.4]
	  assign _T_458 = _T_153 ? 2'h1 : _T_457; // @[Lookup.scala 11:37:@336.4]
	  assign _T_459 = _T_149 ? 2'h1 : _T_458; // @[Lookup.scala 11:37:@337.4]
	  assign _T_460 = _T_145 ? 2'h1 : _T_459; // @[Lookup.scala 11:37:@338.4]
	  assign _T_461 = _T_141 ? 2'h1 : _T_460; // @[Lookup.scala 11:37:@339.4]
	  assign _T_462 = _T_137 ? 2'h1 : _T_461; // @[Lookup.scala 11:37:@340.4]
	  assign _T_463 = _T_133 ? 2'h1 : _T_462; // @[Lookup.scala 11:37:@341.4]
	  assign _T_464 = _T_129 ? 2'h1 : _T_463; // @[Lookup.scala 11:37:@342.4]
	  assign _T_465 = _T_125 ? 2'h1 : _T_464; // @[Lookup.scala 11:37:@343.4]
	  assign _T_466 = _T_121 ? 2'h0 : _T_465; // @[Lookup.scala 11:37:@344.4]
	  assign _T_467 = _T_117 ? 2'h3 : _T_466; // @[Lookup.scala 11:37:@345.4]
	  assign _T_468 = _T_113 ? 2'h2 : _T_467; // @[Lookup.scala 11:37:@346.4]
	  assign _T_469 = _T_109 ? 2'h2 : _T_468; // @[Lookup.scala 11:37:@347.4]
	  assign _T_470 = _T_105 ? 2'h2 : _T_469; // @[Lookup.scala 11:37:@348.4]
	  assign _T_471 = _T_101 ? 2'h1 : _T_470; // @[Lookup.scala 11:37:@349.4]
	  assign _T_472 = _T_97 ? 2'h1 : _T_471; // @[Lookup.scala 11:37:@350.4]
	  assign _T_473 = _T_93 ? 2'h1 : _T_472; // @[Lookup.scala 11:37:@351.4]
	  assign _T_481 = _T_253 ? 4'h8 : 4'h0; // @[Lookup.scala 11:37:@360.4]
	  assign _T_482 = _T_249 ? 4'h8 : _T_481; // @[Lookup.scala 11:37:@361.4]
	  assign _T_483 = _T_245 ? 4'h8 : _T_482; // @[Lookup.scala 11:37:@362.4]
	  assign _T_484 = _T_241 ? 4'h8 : _T_483; // @[Lookup.scala 11:37:@363.4]
	  assign _T_485 = _T_237 ? 4'h8 : _T_484; // @[Lookup.scala 11:37:@364.4]
	  assign _T_486 = _T_233 ? 4'h8 : _T_485; // @[Lookup.scala 11:37:@365.4]
	  assign _T_487 = _T_229 ? 5'h12 : {{1'd0}, _T_486}; // @[Lookup.scala 11:37:@366.4]
	  assign _T_488 = _T_225 ? 5'h11 : _T_487; // @[Lookup.scala 11:37:@367.4]
	  assign _T_489 = _T_221 ? 5'h12 : _T_488; // @[Lookup.scala 11:37:@368.4]
	  assign _T_490 = _T_217 ? 5'h11 : _T_489; // @[Lookup.scala 11:37:@369.4]
	  assign _T_491 = _T_213 ? 5'h10 : _T_490; // @[Lookup.scala 11:37:@370.4]
	  assign _T_492 = _T_209 ? 5'h10 : _T_491; // @[Lookup.scala 11:37:@371.4]
	  assign _T_493 = _T_205 ? 5'h0 : _T_492; // @[Lookup.scala 11:37:@372.4]
	  assign _T_494 = _T_201 ? 5'h0 : _T_493; // @[Lookup.scala 11:37:@373.4]
	  assign _T_495 = _T_197 ? 5'h5 : _T_494; // @[Lookup.scala 11:37:@374.4]
	  assign _T_496 = _T_193 ? 5'h6 : _T_495; // @[Lookup.scala 11:37:@375.4]
	  assign _T_497 = _T_189 ? 5'h1 : _T_496; // @[Lookup.scala 11:37:@376.4]
	  assign _T_498 = _T_185 ? 5'h2 : _T_497; // @[Lookup.scala 11:37:@377.4]
	  assign _T_499 = _T_181 ? 5'h3 : _T_498; // @[Lookup.scala 11:37:@378.4]
	  assign _T_500 = _T_177 ? 5'h12 : _T_499; // @[Lookup.scala 11:37:@379.4]
	  assign _T_501 = _T_173 ? 5'h11 : _T_500; // @[Lookup.scala 11:37:@380.4]
	  assign _T_502 = _T_169 ? 5'h10 : _T_501; // @[Lookup.scala 11:37:@381.4]
	  assign _T_503 = _T_165 ? 5'h0 : _T_502; // @[Lookup.scala 11:37:@382.4]
	  assign _T_504 = _T_161 ? 5'h4 : _T_503; // @[Lookup.scala 11:37:@383.4]
	  assign _T_505 = _T_157 ? 5'h5 : _T_504; // @[Lookup.scala 11:37:@384.4]
	  assign _T_506 = _T_153 ? 5'h6 : _T_505; // @[Lookup.scala 11:37:@385.4]
	  assign _T_507 = _T_149 ? 5'h4 : _T_506; // @[Lookup.scala 11:37:@386.4]
	  assign _T_508 = _T_145 ? 5'h12 : _T_507; // @[Lookup.scala 11:37:@387.4]
	  assign _T_509 = _T_141 ? 5'h11 : _T_508; // @[Lookup.scala 11:37:@388.4]
	  assign _T_510 = _T_137 ? 5'h1 : _T_509; // @[Lookup.scala 11:37:@389.4]
	  assign _T_511 = _T_133 ? 5'h2 : _T_510; // @[Lookup.scala 11:37:@390.4]
	  assign _T_512 = _T_129 ? 5'h3 : _T_511; // @[Lookup.scala 11:37:@391.4]
	  assign _T_513 = _T_125 ? 5'h0 : _T_512; // @[Lookup.scala 11:37:@392.4]
	  assign _T_514 = _T_121 ? 5'h8 : _T_513; // @[Lookup.scala 11:37:@393.4]
	  assign _T_515 = _T_117 ? 5'h0 : _T_514; // @[Lookup.scala 11:37:@394.4]
	  assign _T_516 = _T_113 ? 5'h0 : _T_515; // @[Lookup.scala 11:37:@395.4]
	  assign _T_517 = _T_109 ? 5'h0 : _T_516; // @[Lookup.scala 11:37:@396.4]
	  assign _T_518 = _T_105 ? 5'h0 : _T_517; // @[Lookup.scala 11:37:@397.4]
	  assign _T_519 = _T_101 ? 5'h0 : _T_518; // @[Lookup.scala 11:37:@398.4]
	  assign _T_520 = _T_97 ? 5'h0 : _T_519; // @[Lookup.scala 11:37:@399.4]
	  assign _T_521 = _T_93 ? 5'h0 : _T_520; // @[Lookup.scala 11:37:@400.4]
	  assign csignals_4 = _T_89 ? 5'h0 : _T_521; // @[Lookup.scala 11:37:@401.4]
	  assign _T_529 = _T_253 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@409.4]
	  assign _T_530 = _T_249 ? 2'h3 : _T_529; // @[Lookup.scala 11:37:@410.4]
	  assign _T_531 = _T_245 ? 2'h3 : _T_530; // @[Lookup.scala 11:37:@411.4]
	  assign _T_532 = _T_241 ? 2'h3 : _T_531; // @[Lookup.scala 11:37:@412.4]
	  assign _T_533 = _T_237 ? 2'h3 : _T_532; // @[Lookup.scala 11:37:@413.4]
	  assign _T_534 = _T_233 ? 2'h3 : _T_533; // @[Lookup.scala 11:37:@414.4]
	  assign _T_535 = _T_229 ? 2'h0 : _T_534; // @[Lookup.scala 11:37:@415.4]
	  assign _T_536 = _T_225 ? 2'h0 : _T_535; // @[Lookup.scala 11:37:@416.4]
	  assign _T_537 = _T_221 ? 2'h0 : _T_536; // @[Lookup.scala 11:37:@417.4]
	  assign _T_538 = _T_217 ? 2'h0 : _T_537; // @[Lookup.scala 11:37:@418.4]
	  assign _T_539 = _T_213 ? 2'h0 : _T_538; // @[Lookup.scala 11:37:@419.4]
	  assign _T_540 = _T_209 ? 2'h0 : _T_539; // @[Lookup.scala 11:37:@420.4]
	  assign _T_541 = _T_205 ? 2'h2 : _T_540; // @[Lookup.scala 11:37:@421.4]
	  assign _T_542 = _T_201 ? 2'h2 : _T_541; // @[Lookup.scala 11:37:@422.4]
	  assign _T_543 = _T_197 ? 2'h0 : _T_542; // @[Lookup.scala 11:37:@423.4]
	  assign _T_544 = _T_193 ? 2'h0 : _T_543; // @[Lookup.scala 11:37:@424.4]
	  assign _T_545 = _T_189 ? 2'h0 : _T_544; // @[Lookup.scala 11:37:@425.4]
	  assign _T_546 = _T_185 ? 2'h0 : _T_545; // @[Lookup.scala 11:37:@426.4]
	  assign _T_547 = _T_181 ? 2'h0 : _T_546; // @[Lookup.scala 11:37:@427.4]
	  assign _T_548 = _T_177 ? 2'h0 : _T_547; // @[Lookup.scala 11:37:@428.4]
	  assign _T_549 = _T_173 ? 2'h0 : _T_548; // @[Lookup.scala 11:37:@429.4]
	  assign _T_550 = _T_169 ? 2'h0 : _T_549; // @[Lookup.scala 11:37:@430.4]
	  assign _T_551 = _T_165 ? 2'h0 : _T_550; // @[Lookup.scala 11:37:@431.4]
	  assign _T_552 = _T_161 ? 2'h0 : _T_551; // @[Lookup.scala 11:37:@432.4]
	  assign _T_553 = _T_157 ? 2'h0 : _T_552; // @[Lookup.scala 11:37:@433.4]
	  assign _T_554 = _T_153 ? 2'h0 : _T_553; // @[Lookup.scala 11:37:@434.4]
	  assign _T_555 = _T_149 ? 2'h0 : _T_554; // @[Lookup.scala 11:37:@435.4]
	  assign _T_556 = _T_145 ? 2'h0 : _T_555; // @[Lookup.scala 11:37:@436.4]
	  assign _T_557 = _T_141 ? 2'h0 : _T_556; // @[Lookup.scala 11:37:@437.4]
	  assign _T_558 = _T_137 ? 2'h0 : _T_557; // @[Lookup.scala 11:37:@438.4]
	  assign _T_559 = _T_133 ? 2'h0 : _T_558; // @[Lookup.scala 11:37:@439.4]
	  assign _T_560 = _T_129 ? 2'h0 : _T_559; // @[Lookup.scala 11:37:@440.4]
	  assign _T_561 = _T_125 ? 2'h0 : _T_560; // @[Lookup.scala 11:37:@441.4]
	  assign _T_562 = _T_121 ? 2'h0 : _T_561; // @[Lookup.scala 11:37:@442.4]
	  assign _T_563 = _T_117 ? 2'h0 : _T_562; // @[Lookup.scala 11:37:@443.4]
	  assign _T_564 = _T_113 ? 2'h0 : _T_563; // @[Lookup.scala 11:37:@444.4]
	  assign _T_565 = _T_109 ? 2'h0 : _T_564; // @[Lookup.scala 11:37:@445.4]
	  assign _T_566 = _T_105 ? 2'h0 : _T_565; // @[Lookup.scala 11:37:@446.4]
	  assign _T_567 = _T_101 ? 2'h1 : _T_566; // @[Lookup.scala 11:37:@447.4]
	  assign _T_568 = _T_97 ? 2'h1 : _T_567; // @[Lookup.scala 11:37:@448.4]
	  assign _T_569 = _T_93 ? 2'h1 : _T_568; // @[Lookup.scala 11:37:@449.4]
	  assign _T_578 = _T_249 ? 1'h1 : _T_253; // @[Lookup.scala 11:37:@459.4]
	  assign _T_579 = _T_245 ? 1'h1 : _T_578; // @[Lookup.scala 11:37:@460.4]
	  assign _T_580 = _T_241 ? 1'h1 : _T_579; // @[Lookup.scala 11:37:@461.4]
	  assign _T_581 = _T_237 ? 1'h1 : _T_580; // @[Lookup.scala 11:37:@462.4]
	  assign _T_582 = _T_233 ? 1'h1 : _T_581; // @[Lookup.scala 11:37:@463.4]
	  assign _T_583 = _T_229 ? 1'h0 : _T_582; // @[Lookup.scala 11:37:@464.4]
	  assign _T_584 = _T_225 ? 1'h0 : _T_583; // @[Lookup.scala 11:37:@465.4]
	  assign _T_585 = _T_221 ? 1'h0 : _T_584; // @[Lookup.scala 11:37:@466.4]
	  assign _T_586 = _T_217 ? 1'h0 : _T_585; // @[Lookup.scala 11:37:@467.4]
	  assign _T_587 = _T_213 ? 1'h0 : _T_586; // @[Lookup.scala 11:37:@468.4]
	  assign _T_588 = _T_209 ? 1'h0 : _T_587; // @[Lookup.scala 11:37:@469.4]
	  assign _T_589 = _T_205 ? 1'h1 : _T_588; // @[Lookup.scala 11:37:@470.4]
	  assign _T_590 = _T_201 ? 1'h1 : _T_589; // @[Lookup.scala 11:37:@471.4]
	  assign _T_591 = _T_197 ? 1'h1 : _T_590; // @[Lookup.scala 11:37:@472.4]
	  assign _T_592 = _T_193 ? 1'h1 : _T_591; // @[Lookup.scala 11:37:@473.4]
	  assign _T_593 = _T_189 ? 1'h1 : _T_592; // @[Lookup.scala 11:37:@474.4]
	  assign _T_594 = _T_185 ? 1'h1 : _T_593; // @[Lookup.scala 11:37:@475.4]
	  assign _T_595 = _T_181 ? 1'h1 : _T_594; // @[Lookup.scala 11:37:@476.4]
	  assign _T_596 = _T_177 ? 1'h1 : _T_595; // @[Lookup.scala 11:37:@477.4]
	  assign _T_597 = _T_173 ? 1'h1 : _T_596; // @[Lookup.scala 11:37:@478.4]
	  assign _T_598 = _T_169 ? 1'h1 : _T_597; // @[Lookup.scala 11:37:@479.4]
	  assign _T_599 = _T_165 ? 1'h1 : _T_598; // @[Lookup.scala 11:37:@480.4]
	  assign _T_600 = _T_161 ? 1'h1 : _T_599; // @[Lookup.scala 11:37:@481.4]
	  assign _T_601 = _T_157 ? 1'h1 : _T_600; // @[Lookup.scala 11:37:@482.4]
	  assign _T_602 = _T_153 ? 1'h1 : _T_601; // @[Lookup.scala 11:37:@483.4]
	  assign _T_603 = _T_149 ? 1'h1 : _T_602; // @[Lookup.scala 11:37:@484.4]
	  assign _T_604 = _T_145 ? 1'h1 : _T_603; // @[Lookup.scala 11:37:@485.4]
	  assign _T_605 = _T_141 ? 1'h1 : _T_604; // @[Lookup.scala 11:37:@486.4]
	  assign _T_606 = _T_137 ? 1'h1 : _T_605; // @[Lookup.scala 11:37:@487.4]
	  assign _T_607 = _T_133 ? 1'h1 : _T_606; // @[Lookup.scala 11:37:@488.4]
	  assign _T_608 = _T_129 ? 1'h1 : _T_607; // @[Lookup.scala 11:37:@489.4]
	  assign _T_609 = _T_125 ? 1'h1 : _T_608; // @[Lookup.scala 11:37:@490.4]
	  assign _T_610 = _T_121 ? 1'h1 : _T_609; // @[Lookup.scala 11:37:@491.4]
	  assign _T_611 = _T_117 ? 1'h1 : _T_610; // @[Lookup.scala 11:37:@492.4]
	  assign _T_612 = _T_113 ? 1'h0 : _T_611; // @[Lookup.scala 11:37:@493.4]
	  assign _T_613 = _T_109 ? 1'h0 : _T_612; // @[Lookup.scala 11:37:@494.4]
	  assign _T_614 = _T_105 ? 1'h0 : _T_613; // @[Lookup.scala 11:37:@495.4]
	  assign _T_615 = _T_101 ? 1'h1 : _T_614; // @[Lookup.scala 11:37:@496.4]
	  assign _T_616 = _T_97 ? 1'h1 : _T_615; // @[Lookup.scala 11:37:@497.4]
	  assign _T_617 = _T_93 ? 1'h1 : _T_616; // @[Lookup.scala 11:37:@498.4]
	  assign _T_619 = _T_277 ? 1'h0 : _T_281; // @[Lookup.scala 11:37:@501.4]
	  assign _T_620 = _T_273 ? 1'h0 : _T_619; // @[Lookup.scala 11:37:@502.4]
	  assign _T_621 = _T_269 ? 1'h0 : _T_620; // @[Lookup.scala 11:37:@503.4]
	  assign _T_622 = _T_265 ? 1'h0 : _T_621; // @[Lookup.scala 11:37:@504.4]
	  assign _T_623 = _T_261 ? 1'h0 : _T_622; // @[Lookup.scala 11:37:@505.4]
	  assign _T_624 = _T_257 ? 1'h0 : _T_623; // @[Lookup.scala 11:37:@506.4]
	  assign _T_625 = _T_253 ? 1'h0 : _T_624; // @[Lookup.scala 11:37:@507.4]
	  assign _T_626 = _T_249 ? 1'h0 : _T_625; // @[Lookup.scala 11:37:@508.4]
	  assign _T_627 = _T_245 ? 1'h0 : _T_626; // @[Lookup.scala 11:37:@509.4]
	  assign _T_628 = _T_241 ? 1'h0 : _T_627; // @[Lookup.scala 11:37:@510.4]
	  assign _T_629 = _T_237 ? 1'h0 : _T_628; // @[Lookup.scala 11:37:@511.4]
	  assign _T_630 = _T_233 ? 1'h0 : _T_629; // @[Lookup.scala 11:37:@512.4]
	  assign _T_631 = _T_229 ? 1'h0 : _T_630; // @[Lookup.scala 11:37:@513.4]
	  assign _T_632 = _T_225 ? 1'h0 : _T_631; // @[Lookup.scala 11:37:@514.4]
	  assign _T_633 = _T_221 ? 1'h0 : _T_632; // @[Lookup.scala 11:37:@515.4]
	  assign _T_634 = _T_217 ? 1'h0 : _T_633; // @[Lookup.scala 11:37:@516.4]
	  assign _T_635 = _T_213 ? 1'h0 : _T_634; // @[Lookup.scala 11:37:@517.4]
	  assign _T_636 = _T_209 ? 1'h0 : _T_635; // @[Lookup.scala 11:37:@518.4]
	  assign _T_637 = _T_205 ? 1'h0 : _T_636; // @[Lookup.scala 11:37:@519.4]
	  assign _T_638 = _T_201 ? 1'h0 : _T_637; // @[Lookup.scala 11:37:@520.4]
	  assign _T_639 = _T_197 ? 1'h0 : _T_638; // @[Lookup.scala 11:37:@521.4]
	  assign _T_640 = _T_193 ? 1'h0 : _T_639; // @[Lookup.scala 11:37:@522.4]
	  assign _T_641 = _T_189 ? 1'h0 : _T_640; // @[Lookup.scala 11:37:@523.4]
	  assign _T_642 = _T_185 ? 1'h0 : _T_641; // @[Lookup.scala 11:37:@524.4]
	  assign _T_643 = _T_181 ? 1'h0 : _T_642; // @[Lookup.scala 11:37:@525.4]
	  assign _T_644 = _T_177 ? 1'h0 : _T_643; // @[Lookup.scala 11:37:@526.4]
	  assign _T_645 = _T_173 ? 1'h0 : _T_644; // @[Lookup.scala 11:37:@527.4]
	  assign _T_646 = _T_169 ? 1'h0 : _T_645; // @[Lookup.scala 11:37:@528.4]
	  assign _T_647 = _T_165 ? 1'h0 : _T_646; // @[Lookup.scala 11:37:@529.4]
	  assign _T_648 = _T_161 ? 1'h0 : _T_647; // @[Lookup.scala 11:37:@530.4]
	  assign _T_649 = _T_157 ? 1'h0 : _T_648; // @[Lookup.scala 11:37:@531.4]
	  assign _T_650 = _T_153 ? 1'h0 : _T_649; // @[Lookup.scala 11:37:@532.4]
	  assign _T_651 = _T_149 ? 1'h0 : _T_650; // @[Lookup.scala 11:37:@533.4]
	  assign _T_652 = _T_145 ? 1'h0 : _T_651; // @[Lookup.scala 11:37:@534.4]
	  assign _T_653 = _T_141 ? 1'h0 : _T_652; // @[Lookup.scala 11:37:@535.4]
	  assign _T_654 = _T_137 ? 1'h0 : _T_653; // @[Lookup.scala 11:37:@536.4]
	  assign _T_655 = _T_133 ? 1'h0 : _T_654; // @[Lookup.scala 11:37:@537.4]
	  assign _T_656 = _T_129 ? 1'h0 : _T_655; // @[Lookup.scala 11:37:@538.4]
	  assign _T_657 = _T_125 ? 1'h0 : _T_656; // @[Lookup.scala 11:37:@539.4]
	  assign _T_658 = _T_121 ? 1'h0 : _T_657; // @[Lookup.scala 11:37:@540.4]
	  assign _T_659 = _T_117 ? 1'h0 : _T_658; // @[Lookup.scala 11:37:@541.4]
	  assign _T_660 = _T_113 ? 1'h1 : _T_659; // @[Lookup.scala 11:37:@542.4]
	  assign _T_661 = _T_109 ? 1'h1 : _T_660; // @[Lookup.scala 11:37:@543.4]
	  assign _T_662 = _T_105 ? 1'h1 : _T_661; // @[Lookup.scala 11:37:@544.4]
	  assign _T_663 = _T_101 ? 1'h1 : _T_662; // @[Lookup.scala 11:37:@545.4]
	  assign _T_664 = _T_97 ? 1'h1 : _T_663; // @[Lookup.scala 11:37:@546.4]
	  assign _T_665 = _T_93 ? 1'h1 : _T_664; // @[Lookup.scala 11:37:@547.4]
	  assign _T_709 = _T_109 ? 1'h1 : _T_113; // @[Lookup.scala 11:37:@592.4]
	  assign _T_710 = _T_105 ? 1'h1 : _T_709; // @[Lookup.scala 11:37:@593.4]
	  assign _T_711 = _T_101 ? 1'h0 : _T_710; // @[Lookup.scala 11:37:@594.4]
	  assign _T_712 = _T_97 ? 1'h0 : _T_711; // @[Lookup.scala 11:37:@595.4]
	  assign _T_713 = _T_93 ? 1'h0 : _T_712; // @[Lookup.scala 11:37:@596.4]
	  assign _T_756 = _T_113 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37:@640.4]
	  assign _T_757 = _T_109 ? 3'h1 : _T_756; // @[Lookup.scala 11:37:@641.4]
	  assign _T_758 = _T_105 ? 3'h3 : _T_757; // @[Lookup.scala 11:37:@642.4]
	  assign _T_759 = _T_101 ? 3'h6 : _T_758; // @[Lookup.scala 11:37:@643.4]
	  assign _T_760 = _T_97 ? 3'h5 : _T_759; // @[Lookup.scala 11:37:@644.4]
	  assign _T_761 = _T_93 ? 3'h1 : _T_760; // @[Lookup.scala 11:37:@645.4]
	  assign io_br_type = _T_89 ? 4'h0 : _T_377; // @[IDU.scala 91:21:@697.4]
	  assign io_op1_sel = _T_89 ? 2'h0 : _T_425; // @[IDU.scala 92:21:@698.4]
	  assign io_op2_sel = _T_89 ? 2'h1 : _T_473; // @[IDU.scala 93:21:@699.4]
	  assign io_alu_op = {{1'd0}, csignals_4}; // @[IDU.scala 94:21:@700.4]
	  assign io_wb_sel = _T_89 ? 2'h1 : _T_569; // @[IDU.scala 95:21:@701.4]
	  assign io_rf_wen = _T_89 ? 1'h1 : _T_617; // @[IDU.scala 96:21:@702.4]
	  assign io_mem_en = _T_89 ? 1'h1 : _T_665; // @[IDU.scala 97:21:@703.4]
	  assign io_mem_fcn = _T_89 ? 1'h0 : _T_713; // @[IDU.scala 98:21:@704.4]
	  assign io_mem_msk = _T_89 ? 3'h3 : _T_761; // @[IDU.scala 99:21:@705.4]
	endmodule
	module RegFile( // @[:@708.2]
 000026	  input         clock, // @[:@709.4]
%000002	  input  [4:0]  io_rs1_addr, // @[:@711.4]
%000060	  output [63:0] io_rs1_data, // @[:@711.4]
%000007	  input  [4:0]  io_rs2_addr, // @[:@711.4]
%000000	  output [63:0] io_rs2_data, // @[:@711.4]
%000006	  input  [4:0]  io_waddr, // @[:@711.4]
%000067	  input  [63:0] io_wdata, // @[:@711.4]
%000001	  input         io_wen // @[:@711.4]
	);
	  reg [63:0] regfile [0:31]; // @[RegFile.scala 19:22:@713.4]
	  reg [63:0] _RAND_0;
%000063	  wire [63:0] regfile__T_24_data; // @[RegFile.scala 19:22:@713.4]
%000002	  wire [4:0] regfile__T_24_addr; // @[RegFile.scala 19:22:@713.4]
%000000	  wire [63:0] regfile__T_29_data; // @[RegFile.scala 19:22:@713.4]
%000007	  wire [4:0] regfile__T_29_addr; // @[RegFile.scala 19:22:@713.4]
%000067	  wire [63:0] regfile__T_21_data; // @[RegFile.scala 19:22:@713.4]
%000006	  wire [4:0] regfile__T_21_addr; // @[RegFile.scala 19:22:@713.4]
%000001	  wire  regfile__T_21_mask; // @[RegFile.scala 19:22:@713.4]
%000001	  wire  regfile__T_21_en; // @[RegFile.scala 19:22:@713.4]
	  wire  _T_23; // @[RegFile.scala 22:37:@718.4]
	  wire  _T_28; // @[RegFile.scala 23:37:@722.4]
	  assign regfile__T_24_addr = io_rs1_addr;
	  assign regfile__T_24_data = regfile[regfile__T_24_addr]; // @[RegFile.scala 19:22:@713.4]
	  assign regfile__T_29_addr = io_rs2_addr;
	  assign regfile__T_29_data = regfile[regfile__T_29_addr]; // @[RegFile.scala 19:22:@713.4]
	  assign regfile__T_21_data = io_wdata;
	  assign regfile__T_21_addr = io_waddr;
	  assign regfile__T_21_mask = 1'h1;
	  assign regfile__T_21_en = io_wen;
	  assign _T_23 = io_rs1_addr != 5'h0; // @[RegFile.scala 22:37:@718.4]
	  assign _T_28 = io_rs2_addr != 5'h0; // @[RegFile.scala 23:37:@722.4]
	  assign io_rs1_data = _T_23 ? regfile__T_24_data : 64'h0; // @[RegFile.scala 22:17:@721.4]
	  assign io_rs2_data = _T_28 ? regfile__T_29_data : 64'h0; // @[RegFile.scala 23:17:@725.4]
	`ifdef RANDOMIZE_GARBAGE_ASSIGN
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE_INVALID_ASSIGN
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE_REG_INIT
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE_MEM_INIT
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE
	  integer initvar;
	  initial begin
	    `ifndef verilator
	      #0.002 begin end
	    `endif
	  _RAND_0 = {2{$random}};
	  `ifdef RANDOMIZE_MEM_INIT
	  for (initvar = 0; initvar < 32; initvar = initvar+1)
	    regfile[initvar] = _RAND_0[63:0];
	  `endif // RANDOMIZE_MEM_INIT
	  end
	`endif // RANDOMIZE
 000024	  always @(posedge clock) begin
 000024	    if(regfile__T_21_en & regfile__T_21_mask) begin
%000000	    verilator_coverage: (next point on previous line)

 000012	      regfile[regfile__T_21_addr] <= regfile__T_21_data; // @[RegFile.scala 19:22:@713.4]
	    end
	  end
	endmodule
	module Top( // @[:@727.2]
 000026	  input         clock, // @[:@728.4]
%000002	  input         reset, // @[:@729.4]
%000001	  input         io_imem_req_ready, // @[:@730.4]
%000001	  output        io_imem_req_valid, // @[:@730.4]
%000018	  output [31:0] io_imem_req_bits_addr, // @[:@730.4]
%000000	  output [31:0] io_imem_req_bits_data, // @[:@730.4]
%000000	  output        io_imem_req_bits_fcn, // @[:@730.4]
%000003	  output [2:0]  io_imem_req_bits_msk, // @[:@730.4]
%000001	  output        io_imem_resp_ready, // @[:@730.4]
%000001	  input         io_imem_resp_valid, // @[:@730.4]
%000038	  input  [31:0] io_imem_resp_bits_data, // @[:@730.4]
%000000	  input         io_dmem_req_ready, // @[:@730.4]
%000000	  output        io_dmem_req_valid, // @[:@730.4]
%000060	  output [31:0] io_dmem_req_bits_addr, // @[:@730.4]
%000000	  output [63:0] io_dmem_req_bits_data, // @[:@730.4]
%000000	  output        io_dmem_req_bits_fcn, // @[:@730.4]
%000000	  output [2:0]  io_dmem_req_bits_msk, // @[:@730.4]
%000001	  output        io_dmem_resp_ready, // @[:@730.4]
%000000	  input         io_dmem_resp_valid, // @[:@730.4]
%000000	  input  [63:0] io_dmem_resp_bits_data, // @[:@730.4]
%000001	  output        io_debug_io_wen, // @[:@730.4]
%000006	  output [4:0]  io_debug_io_waddr, // @[:@730.4]
%000067	  output [63:0] io_debug_io_wdata, // @[:@730.4]
%000018	  output [63:0] io_debug_io_PC, // @[:@730.4]
%000002	  output        io_debug_io_stall // @[:@730.4]
	);
%000002	  wire [5:0] alu_io_opcode; // @[core.scala 33:21:@747.4]
%000060	  wire [63:0] alu_io_in1; // @[core.scala 33:21:@747.4]
%000060	  wire [63:0] alu_io_in2; // @[core.scala 33:21:@747.4]
%000062	  wire [63:0] alu_io_out; // @[core.scala 33:21:@747.4]
%000003	  wire  alu_io_zero; // @[core.scala 33:21:@747.4]
%000042	  wire [31:0] idu_io_inst; // @[core.scala 34:21:@750.4]
%000003	  wire [3:0] idu_io_br_type; // @[core.scala 34:21:@750.4]
%000000	  wire [1:0] idu_io_op1_sel; // @[core.scala 34:21:@750.4]
%000002	  wire [1:0] idu_io_op2_sel; // @[core.scala 34:21:@750.4]
%000002	  wire [5:0] idu_io_alu_op; // @[core.scala 34:21:@750.4]
%000001	  wire [1:0] idu_io_wb_sel; // @[core.scala 34:21:@750.4]
%000001	  wire  idu_io_rf_wen; // @[core.scala 34:21:@750.4]
%000000	  wire  idu_io_mem_en; // @[core.scala 34:21:@750.4]
%000000	  wire  idu_io_mem_fcn; // @[core.scala 34:21:@750.4]
%000000	  wire [2:0] idu_io_mem_msk; // @[core.scala 34:21:@750.4]
 000026	  wire  rf_clock; // @[core.scala 35:21:@753.4]
%000002	  wire [4:0] rf_io_rs1_addr; // @[core.scala 35:21:@753.4]
%000060	  wire [63:0] rf_io_rs1_data; // @[core.scala 35:21:@753.4]
%000007	  wire [4:0] rf_io_rs2_addr; // @[core.scala 35:21:@753.4]
%000000	  wire [63:0] rf_io_rs2_data; // @[core.scala 35:21:@753.4]
%000006	  wire [4:0] rf_io_waddr; // @[core.scala 35:21:@753.4]
%000067	  wire [63:0] rf_io_wdata; // @[core.scala 35:21:@753.4]
%000001	  wire  rf_io_wen; // @[core.scala 35:21:@753.4]
%000018	  reg [63:0] pc_reg; // @[core.scala 17:26:@732.4]
	  reg [63:0] _RAND_0;
	  wire [64:0] _T_100; // @[core.scala 20:23:@735.4]
	  wire [63:0] _T_101; // @[core.scala 20:23:@736.4]
%000042	  wire [31:0] inst; // @[core.scala 29:15:@744.4]
	  wire  _T_108; // @[core.scala 39:17:@757.4]
	  wire  _T_109; // @[core.scala 39:58:@758.4]
	  wire  _T_111; // @[core.scala 39:84:@759.4]
	  wire  _T_112; // @[core.scala 39:81:@760.4]
	  wire  _T_114; // @[core.scala 39:40:@761.4]
%000002	  wire  stall; // @[core.scala 39:37:@762.4]
%000022	  wire [11:0] imm_i; // @[core.scala 42:21:@763.4]
	  wire [6:0] _T_115; // @[core.scala 43:25:@764.4]
	  wire [4:0] _T_116; // @[core.scala 43:39:@765.4]
%000021	  wire [11:0] imm_s; // @[Cat.scala 30:58:@766.4]
	  wire  _T_117; // @[core.scala 44:25:@767.4]
	  wire  _T_118; // @[core.scala 44:35:@768.4]
	  wire [5:0] _T_119; // @[core.scala 44:44:@769.4]
	  wire [3:0] _T_120; // @[core.scala 44:57:@770.4]
	  wire [9:0] _T_121; // @[Cat.scala 30:58:@771.4]
	  wire [1:0] _T_122; // @[Cat.scala 30:58:@772.4]
%000021	  wire [11:0] imm_b; // @[Cat.scala 30:58:@773.4]
%000026	  wire [19:0] imm_u; // @[core.scala 45:21:@774.4]
	  wire [7:0] _T_124; // @[core.scala 46:35:@776.4]
	  wire  _T_125; // @[core.scala 46:48:@777.4]
	  wire [9:0] _T_126; // @[core.scala 46:58:@778.4]
	  wire [10:0] _T_127; // @[Cat.scala 30:58:@779.4]
	  wire [8:0] _T_128; // @[Cat.scala 30:58:@780.4]
%000026	  wire [19:0] imm_j; // @[Cat.scala 30:58:@781.4]
	  wire [4:0] _T_134; // @[core.scala 47:39:@783.4]
%000002	  wire [31:0] imm_z; // @[Cat.scala 30:58:@784.4]
	  wire  _T_135; // @[core.scala 50:39:@785.4]
	  wire [19:0] _T_139; // @[Bitwise.scala 72:12:@787.4]
%000062	  wire [31:0] imm_i_sext; // @[Cat.scala 30:58:@788.4]
	  wire  _T_140; // @[core.scala 51:39:@789.4]
	  wire [19:0] _T_144; // @[Bitwise.scala 72:12:@791.4]
%000061	  wire [31:0] imm_s_sext; // @[Cat.scala 30:58:@792.4]
	  wire  _T_145; // @[core.scala 52:39:@793.4]
	  wire [18:0] _T_149; // @[Bitwise.scala 72:12:@795.4]
	  wire [30:0] _T_151; // @[Cat.scala 30:58:@796.4]
%000059	  wire [31:0] imm_b_sext; // @[Cat.scala 30:58:@797.4]
%000026	  wire [31:0] imm_u_sext; // @[Cat.scala 30:58:@799.4]
	  wire  _T_157; // @[core.scala 54:39:@800.4]
	  wire [10:0] _T_161; // @[Bitwise.scala 72:12:@802.4]
	  wire [30:0] _T_163; // @[Cat.scala 30:58:@803.4]
%000048	  wire [31:0] imm_j_sext; // @[Cat.scala 30:58:@804.4]
	  wire  _T_167; // @[core.scala 61:24:@811.4]
	  wire  _T_168; // @[core.scala 62:24:@812.4]
	  wire  _T_169; // @[core.scala 63:24:@813.4]
%000019	  wire [31:0] pc_4; // @[core.scala 19:23:@734.4 core.scala 20:13:@737.4]
	  wire [63:0] _T_170; // @[Mux.scala 61:16:@814.4]
	  wire [63:0] _T_171; // @[Mux.scala 61:16:@815.4]
	  wire  _T_173; // @[core.scala 70:25:@820.4]
	  wire  _T_174; // @[core.scala 71:25:@821.4]
	  wire  _T_175; // @[core.scala 72:25:@822.4]
	  wire [63:0] _T_176; // @[Mux.scala 61:16:@823.4]
	  wire [63:0] _T_177; // @[Mux.scala 61:16:@824.4]
	  wire  _T_179; // @[core.scala 76:25:@827.4]
	  wire  _T_180; // @[core.scala 77:25:@828.4]
	  wire  _T_181; // @[core.scala 78:25:@829.4]
	  wire  _T_182; // @[core.scala 79:25:@830.4]
	  wire [63:0] _T_183; // @[Mux.scala 61:16:@831.4]
	  wire [63:0] _T_184; // @[Mux.scala 61:16:@832.4]
	  wire [63:0] _T_185; // @[Mux.scala 61:16:@833.4]
	  wire [63:0] _GEN_1; // @[core.scala 92:29:@842.4]
	  wire [64:0] _T_188; // @[core.scala 92:29:@842.4]
%000072	  wire [63:0] br_target; // @[core.scala 92:29:@843.4]
	  wire [63:0] _GEN_2; // @[core.scala 93:29:@844.4]
	  wire [64:0] _T_189; // @[core.scala 93:29:@844.4]
%000050	  wire [63:0] jmp_target; // @[core.scala 93:29:@845.4]
	  wire [63:0] _GEN_3; // @[core.scala 94:37:@846.4]
	  wire [64:0] _T_190; // @[core.scala 94:37:@846.4]
%000064	  wire [63:0] jr_target; // @[core.scala 94:37:@847.4]
	  wire  _T_192; // @[core.scala 97:25:@848.4]
	  wire  _T_193; // @[core.scala 97:36:@849.4]
	  wire  _T_195; // @[core.scala 98:25:@850.4]
	  wire  _T_197; // @[core.scala 98:39:@851.4]
	  wire  _T_198; // @[core.scala 98:36:@852.4]
	  wire  _T_200; // @[core.scala 99:25:@853.4]
	  wire  _T_201; // @[core.scala 99:50:@854.4]
	  wire  _T_203; // @[core.scala 99:39:@855.4]
	  wire  _T_204; // @[core.scala 99:36:@856.4]
	  wire  _T_206; // @[core.scala 100:25:@857.4]
	  wire  _T_210; // @[core.scala 100:36:@860.4]
	  wire  _T_212; // @[core.scala 101:25:@861.4]
	  wire  _T_214; // @[core.scala 101:36:@863.4]
	  wire  _T_216; // @[core.scala 102:25:@864.4]
	  wire  _T_218; // @[core.scala 102:36:@866.4]
	  wire  _T_221; // @[Mux.scala 61:16:@868.4]
	  wire  _T_222; // @[Mux.scala 61:16:@869.4]
	  wire  _T_223; // @[Mux.scala 61:16:@870.4]
	  wire  _T_224; // @[Mux.scala 61:16:@871.4]
%000000	  wire  br_taken; // @[Mux.scala 61:16:@872.4]
	  wire  _T_227; // @[core.scala 108:25:@874.4]
	  wire  _T_228; // @[core.scala 109:25:@875.4]
	  wire [63:0] _T_229; // @[Mux.scala 61:16:@876.4]
	  wire [63:0] _T_230; // @[Mux.scala 61:16:@877.4]
	  wire [63:0] _T_231; // @[Mux.scala 61:16:@878.4]
	  wire  _T_233; // @[core.scala 111:10:@880.4]
%000022	  wire [31:0] pc_next; // @[core.scala 18:23:@733.4 core.scala 106:13:@879.4]
	  wire [63:0] _GEN_0; // @[core.scala 111:17:@881.4]
	  ALU alu ( // @[core.scala 33:21:@747.4]
	    .io_opcode(alu_io_opcode),
	    .io_in1(alu_io_in1),
	    .io_in2(alu_io_in2),
	    .io_out(alu_io_out),
	    .io_zero(alu_io_zero)
	  );
	  IDU idu ( // @[core.scala 34:21:@750.4]
	    .io_inst(idu_io_inst),
	    .io_br_type(idu_io_br_type),
	    .io_op1_sel(idu_io_op1_sel),
	    .io_op2_sel(idu_io_op2_sel),
	    .io_alu_op(idu_io_alu_op),
	    .io_wb_sel(idu_io_wb_sel),
	    .io_rf_wen(idu_io_rf_wen),
	    .io_mem_en(idu_io_mem_en),
	    .io_mem_fcn(idu_io_mem_fcn),
	    .io_mem_msk(idu_io_mem_msk)
	  );
	  RegFile rf ( // @[core.scala 35:21:@753.4]
	    .clock(rf_clock),
	    .io_rs1_addr(rf_io_rs1_addr),
	    .io_rs1_data(rf_io_rs1_data),
	    .io_rs2_addr(rf_io_rs2_addr),
	    .io_rs2_data(rf_io_rs2_data),
	    .io_waddr(rf_io_waddr),
	    .io_wdata(rf_io_wdata),
	    .io_wen(rf_io_wen)
	  );
	  assign _T_100 = pc_reg + 64'h4; // @[core.scala 20:23:@735.4]
	  assign _T_101 = _T_100[63:0]; // @[core.scala 20:23:@736.4]
	  assign inst = io_imem_resp_valid ? io_imem_resp_bits_data : 32'h4033; // @[core.scala 29:15:@744.4]
	  assign _T_108 = io_imem_resp_valid == 1'h0; // @[core.scala 39:17:@757.4]
	  assign _T_109 = idu_io_mem_en & io_dmem_resp_valid; // @[core.scala 39:58:@758.4]
	  assign _T_111 = idu_io_mem_en == 1'h0; // @[core.scala 39:84:@759.4]
	  assign _T_112 = _T_109 | _T_111; // @[core.scala 39:81:@760.4]
	  assign _T_114 = _T_112 == 1'h0; // @[core.scala 39:40:@761.4]
	  assign stall = _T_108 | _T_114; // @[core.scala 39:37:@762.4]
	  assign imm_i = inst[31:20]; // @[core.scala 42:21:@763.4]
	  assign _T_115 = inst[31:25]; // @[core.scala 43:25:@764.4]
	  assign _T_116 = inst[11:7]; // @[core.scala 43:39:@765.4]
	  assign imm_s = {_T_115,_T_116}; // @[Cat.scala 30:58:@766.4]
	  assign _T_117 = inst[31]; // @[core.scala 44:25:@767.4]
	  assign _T_118 = inst[7]; // @[core.scala 44:35:@768.4]
	  assign _T_119 = inst[30:25]; // @[core.scala 44:44:@769.4]
	  assign _T_120 = inst[11:8]; // @[core.scala 44:57:@770.4]
	  assign _T_121 = {_T_119,_T_120}; // @[Cat.scala 30:58:@771.4]
	  assign _T_122 = {_T_117,_T_118}; // @[Cat.scala 30:58:@772.4]
	  assign imm_b = {_T_122,_T_121}; // @[Cat.scala 30:58:@773.4]
	  assign imm_u = inst[31:12]; // @[core.scala 45:21:@774.4]
	  assign _T_124 = inst[19:12]; // @[core.scala 46:35:@776.4]
	  assign _T_125 = inst[20]; // @[core.scala 46:48:@777.4]
	  assign _T_126 = inst[30:21]; // @[core.scala 46:58:@778.4]
	  assign _T_127 = {_T_125,_T_126}; // @[Cat.scala 30:58:@779.4]
	  assign _T_128 = {_T_117,_T_124}; // @[Cat.scala 30:58:@780.4]
	  assign imm_j = {_T_128,_T_127}; // @[Cat.scala 30:58:@781.4]
	  assign _T_134 = inst[19:15]; // @[core.scala 47:39:@783.4]
	  assign imm_z = {27'h0,_T_134}; // @[Cat.scala 30:58:@784.4]
	  assign _T_135 = imm_i[11]; // @[core.scala 50:39:@785.4]
	  assign _T_139 = _T_135 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@787.4]
	  assign imm_i_sext = {_T_139,imm_i}; // @[Cat.scala 30:58:@788.4]
	  assign _T_140 = imm_s[11]; // @[core.scala 51:39:@789.4]
	  assign _T_144 = _T_140 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@791.4]
	  assign imm_s_sext = {_T_144,imm_s}; // @[Cat.scala 30:58:@792.4]
	  assign _T_145 = imm_b[11]; // @[core.scala 52:39:@793.4]
	  assign _T_149 = _T_145 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:@795.4]
	  assign _T_151 = {_T_149,imm_b}; // @[Cat.scala 30:58:@796.4]
	  assign imm_b_sext = {_T_151,1'h0}; // @[Cat.scala 30:58:@797.4]
	  assign imm_u_sext = {imm_u,12'h0}; // @[Cat.scala 30:58:@799.4]
	  assign _T_157 = imm_j[19]; // @[core.scala 54:39:@800.4]
	  assign _T_161 = _T_157 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:@802.4]
	  assign _T_163 = {_T_161,imm_j}; // @[Cat.scala 30:58:@803.4]
	  assign imm_j_sext = {_T_163,1'h0}; // @[Cat.scala 30:58:@804.4]
	  assign _T_167 = idu_io_wb_sel == 2'h0; // @[core.scala 61:24:@811.4]
	  assign _T_168 = idu_io_wb_sel == 2'h1; // @[core.scala 62:24:@812.4]
	  assign _T_169 = idu_io_wb_sel == 2'h2; // @[core.scala 63:24:@813.4]
	  assign pc_4 = _T_101[31:0]; // @[core.scala 19:23:@734.4 core.scala 20:13:@737.4]
	  assign _T_170 = _T_169 ? {{32'd0}, pc_4} : alu_io_out; // @[Mux.scala 61:16:@814.4]
	  assign _T_171 = _T_168 ? io_dmem_resp_bits_data : _T_170; // @[Mux.scala 61:16:@815.4]
	  assign _T_173 = idu_io_op1_sel == 2'h0; // @[core.scala 70:25:@820.4]
	  assign _T_174 = idu_io_op1_sel == 2'h1; // @[core.scala 71:25:@821.4]
	  assign _T_175 = idu_io_op1_sel == 2'h2; // @[core.scala 72:25:@822.4]
	  assign _T_176 = _T_175 ? {{32'd0}, imm_z} : rf_io_rs1_data; // @[Mux.scala 61:16:@823.4]
	  assign _T_177 = _T_174 ? {{32'd0}, imm_u_sext} : _T_176; // @[Mux.scala 61:16:@824.4]
	  assign _T_179 = idu_io_op2_sel == 2'h0; // @[core.scala 76:25:@827.4]
	  assign _T_180 = idu_io_op2_sel == 2'h1; // @[core.scala 77:25:@828.4]
	  assign _T_181 = idu_io_op2_sel == 2'h2; // @[core.scala 78:25:@829.4]
	  assign _T_182 = idu_io_op2_sel == 2'h3; // @[core.scala 79:25:@830.4]
	  assign _T_183 = _T_182 ? pc_reg : rf_io_rs2_data; // @[Mux.scala 61:16:@831.4]
	  assign _T_184 = _T_181 ? {{32'd0}, imm_s_sext} : _T_183; // @[Mux.scala 61:16:@832.4]
	  assign _T_185 = _T_180 ? {{32'd0}, imm_i_sext} : _T_184; // @[Mux.scala 61:16:@833.4]
	  assign _GEN_1 = {{32'd0}, imm_b_sext}; // @[core.scala 92:29:@842.4]
	  assign _T_188 = pc_reg + _GEN_1; // @[core.scala 92:29:@842.4]
	  assign br_target = _T_188[63:0]; // @[core.scala 92:29:@843.4]
	  assign _GEN_2 = {{32'd0}, imm_j_sext}; // @[core.scala 93:29:@844.4]
	  assign _T_189 = pc_reg + _GEN_2; // @[core.scala 93:29:@844.4]
	  assign jmp_target = _T_189[63:0]; // @[core.scala 93:29:@845.4]
	  assign _GEN_3 = {{32'd0}, imm_i_sext}; // @[core.scala 94:37:@846.4]
	  assign _T_190 = rf_io_rs1_data + _GEN_3; // @[core.scala 94:37:@846.4]
	  assign jr_target = _T_190[63:0]; // @[core.scala 94:37:@847.4]
	  assign _T_192 = idu_io_br_type == 4'h2; // @[core.scala 97:25:@848.4]
	  assign _T_193 = _T_192 & alu_io_zero; // @[core.scala 97:36:@849.4]
	  assign _T_195 = idu_io_br_type == 4'h1; // @[core.scala 98:25:@850.4]
	  assign _T_197 = alu_io_zero == 1'h0; // @[core.scala 98:39:@851.4]
	  assign _T_198 = _T_195 & _T_197; // @[core.scala 98:36:@852.4]
	  assign _T_200 = idu_io_br_type == 4'h3; // @[core.scala 99:25:@853.4]
	  assign _T_201 = alu_io_out[0]; // @[core.scala 99:50:@854.4]
	  assign _T_203 = _T_201 == 1'h0; // @[core.scala 99:39:@855.4]
	  assign _T_204 = _T_200 & _T_203; // @[core.scala 99:36:@856.4]
	  assign _T_206 = idu_io_br_type == 4'h4; // @[core.scala 100:25:@857.4]
	  assign _T_210 = _T_206 & _T_203; // @[core.scala 100:36:@860.4]
	  assign _T_212 = idu_io_br_type == 4'h5; // @[core.scala 101:25:@861.4]
	  assign _T_214 = _T_212 & _T_201; // @[core.scala 101:36:@863.4]
	  assign _T_216 = idu_io_br_type == 4'h6; // @[core.scala 102:25:@864.4]
	  assign _T_218 = _T_216 & _T_201; // @[core.scala 102:36:@866.4]
	  assign _T_221 = _T_214 ? 1'h1 : _T_218; // @[Mux.scala 61:16:@868.4]
	  assign _T_222 = _T_210 ? 1'h1 : _T_221; // @[Mux.scala 61:16:@869.4]
	  assign _T_223 = _T_204 ? 1'h1 : _T_222; // @[Mux.scala 61:16:@870.4]
	  assign _T_224 = _T_198 ? 1'h1 : _T_223; // @[Mux.scala 61:16:@871.4]
	  assign br_taken = _T_193 ? 1'h1 : _T_224; // @[Mux.scala 61:16:@872.4]
	  assign _T_227 = idu_io_br_type == 4'h7; // @[core.scala 108:25:@874.4]
	  assign _T_228 = idu_io_br_type == 4'h8; // @[core.scala 109:25:@875.4]
	  assign _T_229 = _T_228 ? jr_target : {{32'd0}, pc_4}; // @[Mux.scala 61:16:@876.4]
	  assign _T_230 = _T_227 ? jmp_target : _T_229; // @[Mux.scala 61:16:@877.4]
	  assign _T_231 = br_taken ? br_target : _T_230; // @[Mux.scala 61:16:@878.4]
	  assign _T_233 = stall == 1'h0; // @[core.scala 111:10:@880.4]
	  assign pc_next = _T_231[31:0]; // @[core.scala 18:23:@733.4 core.scala 106:13:@879.4]
	  assign _GEN_0 = _T_233 ? {{32'd0}, pc_next} : pc_reg; // @[core.scala 111:17:@881.4]
	  assign io_imem_req_valid = 1'h1; // @[core.scala 27:29:@742.4]
	  assign io_imem_req_bits_addr = pc_reg[31:0]; // @[core.scala 24:29:@739.4]
	  assign io_imem_req_bits_data = 32'h0; // @[core.scala 23:29:@738.4]
	  assign io_imem_req_bits_fcn = 1'h0; // @[core.scala 25:29:@740.4]
	  assign io_imem_req_bits_msk = 3'h7; // @[core.scala 26:29:@741.4]
	  assign io_imem_resp_ready = 1'h1; // @[core.scala 31:24:@746.4]
	  assign io_dmem_req_valid = idu_io_mem_en; // @[core.scala 85:27:@838.4]
	  assign io_dmem_req_bits_addr = alu_io_out[31:0]; // @[core.scala 83:27:@836.4]
	  assign io_dmem_req_bits_data = rf_io_rs2_data; // @[core.scala 84:27:@837.4]
	  assign io_dmem_req_bits_fcn = idu_io_mem_fcn; // @[core.scala 86:27:@839.4]
	  assign io_dmem_req_bits_msk = idu_io_mem_msk; // @[core.scala 87:27:@840.4]
	  assign io_dmem_resp_ready = 1'h1; // @[core.scala 89:24:@841.4]
	  assign io_debug_io_wen = rf_io_wen; // @[core.scala 116:25:@884.4]
	  assign io_debug_io_waddr = rf_io_waddr; // @[core.scala 117:25:@885.4]
	  assign io_debug_io_wdata = rf_io_wdata; // @[core.scala 118:25:@886.4]
	  assign io_debug_io_PC = pc_reg; // @[core.scala 119:25:@887.4]
	  assign io_debug_io_stall = _T_108 | _T_114; // @[core.scala 120:25:@888.4]
	  assign alu_io_opcode = idu_io_alu_op; // @[core.scala 68:20:@819.4]
	  assign alu_io_in1 = _T_173 ? rf_io_rs1_data : _T_177; // @[core.scala 69:20:@826.4]
	  assign alu_io_in2 = _T_179 ? rf_io_rs2_data : _T_185; // @[core.scala 75:20:@835.4]
	  assign idu_io_inst = io_imem_resp_valid ? io_imem_resp_bits_data : 32'h4033; // @[core.scala 36:17:@756.4]
	  assign rf_clock = clock; // @[:@754.4]
	  assign rf_io_rs1_addr = inst[19:15]; // @[core.scala 57:20:@806.4]
	  assign rf_io_rs2_addr = inst[24:20]; // @[core.scala 58:20:@808.4]
	  assign rf_io_waddr = inst[11:7]; // @[core.scala 59:20:@810.4]
	  assign rf_io_wdata = _T_167 ? alu_io_out : _T_171; // @[core.scala 60:20:@817.4]
	  assign rf_io_wen = idu_io_rf_wen; // @[core.scala 65:20:@818.4]
	`ifdef RANDOMIZE_GARBAGE_ASSIGN
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE_INVALID_ASSIGN
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE_REG_INIT
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE_MEM_INIT
	`define RANDOMIZE
	`endif
	`ifdef RANDOMIZE
	  integer initvar;
	  initial begin
	    `ifndef verilator
	      #0.002 begin end
	    `endif
	  `ifdef RANDOMIZE_REG_INIT
	  _RAND_0 = {2{$random}};
	  pc_reg = _RAND_0[63:0];
	  `endif // RANDOMIZE_REG_INIT
	  end
	`endif // RANDOMIZE
 000024	  always @(posedge clock) begin
%000004	    if (reset) begin
 000010	    verilator_coverage: (next point on previous line)

%000002	      pc_reg <= 64'h80000000;
 000010	    end else begin
%000018	      if (_T_233) begin
%000001	      verilator_coverage: (next point on previous line)

%000009	        pc_reg <= {{32'd0}, pc_next};
	      end
	    end
	  end
%000002	   initial begin
%000002	      if ($test$plusargs("trace") != 0) begin
%000000	      verilator_coverage: (next point on previous line)

%000001	         $display("[%0t] Tracing to logs/vlt_dump.vcd...\n", $time);
%000001	         $dumpfile("logs/vlt_dump.vcd");
%000001	         $dumpvars();
	      end
%000001	      $display("[%0t] Model running...\n", $time);
	   end
	endmodule
	
